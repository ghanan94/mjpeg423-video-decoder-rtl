// ECE423_QSYS.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module ECE423_QSYS (
		input  wire        clk_125_clk,                                  //             clk_125.clk
		input  wire        clk_50_clk,                                   //              clk_50.clk
		output wire        i2c_scl_export,                               //             i2c_scl.export
		inout  wire        i2c_sda_export,                               //             i2c_sda.export
		input  wire [3:0]  key_export,                                   //                 key.export
		output wire [7:0]  ledg_export,                                  //                ledg.export
		output wire [7:0]  ledr_export,                                  //                ledr.export
		output wire [9:0]  lpddr2_mem_ca,                                //              lpddr2.mem_ca
		output wire [0:0]  lpddr2_mem_ck,                                //                    .mem_ck
		output wire [0:0]  lpddr2_mem_ck_n,                              //                    .mem_ck_n
		output wire [0:0]  lpddr2_mem_cke,                               //                    .mem_cke
		output wire [0:0]  lpddr2_mem_cs_n,                              //                    .mem_cs_n
		output wire [3:0]  lpddr2_mem_dm,                                //                    .mem_dm
		inout  wire [31:0] lpddr2_mem_dq,                                //                    .mem_dq
		inout  wire [3:0]  lpddr2_mem_dqs,                               //                    .mem_dqs
		inout  wire [3:0]  lpddr2_mem_dqs_n,                             //                    .mem_dqs_n
		input  wire        lpddr2_global_reset_reset_n,                  // lpddr2_global_reset.reset_n
		input  wire        lpddr2_oct_rzqin,                             //          lpddr2_oct.rzqin
		input  wire        lpddr2_pll_ref_clk_clk,                       //  lpddr2_pll_ref_clk.clk
		output wire        lpddr2_pll_sharing_pll_mem_clk,               //  lpddr2_pll_sharing.pll_mem_clk
		output wire        lpddr2_pll_sharing_pll_write_clk,             //                    .pll_write_clk
		output wire        lpddr2_pll_sharing_pll_locked,                //                    .pll_locked
		output wire        lpddr2_pll_sharing_pll_write_clk_pre_phy_clk, //                    .pll_write_clk_pre_phy_clk
		output wire        lpddr2_pll_sharing_pll_addr_cmd_clk,          //                    .pll_addr_cmd_clk
		output wire        lpddr2_pll_sharing_pll_avl_clk,               //                    .pll_avl_clk
		output wire        lpddr2_pll_sharing_pll_config_clk,            //                    .pll_config_clk
		output wire        lpddr2_pll_sharing_pll_mem_phy_clk,           //                    .pll_mem_phy_clk
		output wire        lpddr2_pll_sharing_afi_phy_clk,               //                    .afi_phy_clk
		output wire        lpddr2_pll_sharing_pll_avl_phy_clk,           //                    .pll_avl_phy_clk
		output wire        lpddr2_status_local_init_done,                //       lpddr2_status.local_init_done
		output wire        lpddr2_status_local_cal_success,              //                    .local_cal_success
		output wire        lpddr2_status_local_cal_fail,                 //                    .local_cal_fail
		input  wire        reset_reset_n,                                //               reset.reset_n
		output wire        sd_sd_clk,                                    //                  sd.sd_clk
		inout  wire        sd_sd_cmd,                                    //                    .sd_cmd
		inout  wire [3:0]  sd_sd_dat,                                    //                    .sd_dat
		inout  wire [15:0] sram_bridge_out_sram_tcm_data_out,            //     sram_bridge_out.sram_tcm_data_out
		output wire [18:0] sram_bridge_out_sram_tcm_address_out,         //                    .sram_tcm_address_out
		output wire [0:0]  sram_bridge_out_sram_tcm_outputenable_n_out,  //                    .sram_tcm_outputenable_n_out
		output wire [0:0]  sram_bridge_out_sram_tcm_chipselect_n_out,    //                    .sram_tcm_chipselect_n_out
		output wire [1:0]  sram_bridge_out_sram_tcm_byteenable_n_out,    //                    .sram_tcm_byteenable_n_out
		output wire [0:0]  sram_bridge_out_sram_tcm_write_n_out,         //                    .sram_tcm_write_n_out
		output wire [23:0] video_RGB_OUT,                                //               video.RGB_OUT
		output wire        video_HD,                                     //                    .HD
		output wire        video_VD,                                     //                    .VD
		output wire        video_DEN,                                    //                    .DEN
		output wire        video_clk_clk                                 //           video_clk.clk
	);

	wire          idct_accelerator_2d_avalon_streaming_source_valid;                            // idct_accelerator_2d:o_valid -> mdma_from_idct_accel:st_sink_valid
	wire   [31:0] idct_accelerator_2d_avalon_streaming_source_data;                             // idct_accelerator_2d:o_data -> mdma_from_idct_accel:st_sink_data
	wire          idct_accelerator_2d_avalon_streaming_source_ready;                            // mdma_from_idct_accel:st_sink_ready -> idct_accelerator_2d:i_ready
	wire          ycbcr_to_rgb_accelerator_avalon_streaming_source_valid;                       // ycbcr_to_rgb_accelerator:o_rgb_valid -> mdma_from_ycbcr_to_rgb_accel:st_sink_valid
	wire   [31:0] ycbcr_to_rgb_accelerator_avalon_streaming_source_data;                        // ycbcr_to_rgb_accelerator:o_rgb_data -> mdma_from_ycbcr_to_rgb_accel:st_sink_data
	wire          ycbcr_to_rgb_accelerator_avalon_streaming_source_ready;                       // mdma_from_ycbcr_to_rgb_accel:st_sink_ready -> ycbcr_to_rgb_accelerator:i_rgb_ready
	wire          pixel_conv_out_valid;                                                         // pixel_conv:valid_out -> video:valid
	wire   [23:0] pixel_conv_out_data;                                                          // pixel_conv:data_out -> video:data
	wire          pixel_conv_out_ready;                                                         // video:ready -> pixel_conv:ready_in
	wire          pixel_conv_out_startofpacket;                                                 // pixel_conv:sop_out -> video:sop
	wire          pixel_conv_out_endofpacket;                                                   // pixel_conv:eop_out -> video:eop
	wire          pixel_conv_out_empty;                                                         // pixel_conv:empty_out -> video:empty
	wire          mdma_to_idct_accel_st_source_valid;                                           // mdma_to_idct_accel:st_source_valid -> idct_accelerator_2d:i_valid
	wire   [31:0] mdma_to_idct_accel_st_source_data;                                            // mdma_to_idct_accel:st_source_data -> idct_accelerator_2d:i_data
	wire          mdma_to_idct_accel_st_source_ready;                                           // idct_accelerator_2d:o_ready -> mdma_to_idct_accel:st_source_ready
	wire          mdma_to_ycbcr_to_rgb_accel_cb_st_source_valid;                                // mdma_to_ycbcr_to_rgb_accel_cb:st_source_valid -> ycbcr_to_rgb_accelerator:i_cb_valid
	wire   [31:0] mdma_to_ycbcr_to_rgb_accel_cb_st_source_data;                                 // mdma_to_ycbcr_to_rgb_accel_cb:st_source_data -> ycbcr_to_rgb_accelerator:i_cb_data
	wire          mdma_to_ycbcr_to_rgb_accel_cb_st_source_ready;                                // ycbcr_to_rgb_accelerator:o_cb_ready -> mdma_to_ycbcr_to_rgb_accel_cb:st_source_ready
	wire          mdma_to_ycbcr_to_rgb_accel_cr_st_source_valid;                                // mdma_to_ycbcr_to_rgb_accel_cr:st_source_valid -> ycbcr_to_rgb_accelerator:i_cr_valid
	wire   [31:0] mdma_to_ycbcr_to_rgb_accel_cr_st_source_data;                                 // mdma_to_ycbcr_to_rgb_accel_cr:st_source_data -> ycbcr_to_rgb_accelerator:i_cr_data
	wire          mdma_to_ycbcr_to_rgb_accel_cr_st_source_ready;                                // ycbcr_to_rgb_accelerator:o_cr_ready -> mdma_to_ycbcr_to_rgb_accel_cr:st_source_ready
	wire          mdma_to_ycbcr_to_rgb_accel_y_st_source_valid;                                 // mdma_to_ycbcr_to_rgb_accel_y:st_source_valid -> ycbcr_to_rgb_accelerator:i_y_valid
	wire   [31:0] mdma_to_ycbcr_to_rgb_accel_y_st_source_data;                                  // mdma_to_ycbcr_to_rgb_accel_y:st_source_data -> ycbcr_to_rgb_accelerator:i_y_data
	wire          mdma_to_ycbcr_to_rgb_accel_y_st_source_ready;                                 // ycbcr_to_rgb_accelerator:o_y_ready -> mdma_to_ycbcr_to_rgb_accel_y:st_source_ready
	wire          reset_controller_0_reset_out_reset;                                           // reset_controller_0:reset_out -> [avalon_st_adapter_001:in_rst_0_reset, i2c_scl:reset_n, i2c_sda:reset_n, idct_accelerator_2d:reset_n, key:reset_n, ledg:reset_n, ledr:reset_n, lpddr2:mp_cmd_reset_n_0_reset_n, lpddr2:mp_cmd_reset_n_1_reset_n, lpddr2:mp_cmd_reset_n_2_reset_n, lpddr2:mp_rfifo_reset_n_0_reset_n, lpddr2:mp_rfifo_reset_n_1_reset_n, lpddr2:mp_wfifo_reset_n_0_reset_n, lpddr2:mp_wfifo_reset_n_1_reset_n, lpddr2:soft_reset_n, mailbox_simple_cpu0_to_cpu1:rst_n, mailbox_simple_cpu1_to_cpu0:rst_n, mdma_from_idct_accel:reset_n_reset_n, mdma_from_ycbcr_to_rgb_accel:reset_n_reset_n, mdma_to_idct_accel:reset_n_reset_n, mdma_to_ycbcr_to_rgb_accel_cb:reset_n_reset_n, mdma_to_ycbcr_to_rgb_accel_cr:reset_n_reset_n, mdma_to_ycbcr_to_rgb_accel_y:reset_n_reset_n, mm_interconnect_0:lpddr2_mp_cmd_reset_n_0_reset_bridge_in_reset_reset, mm_interconnect_0:mailbox_simple_cpu1_to_cpu0_rst_n_reset_bridge_in_reset_reset, mm_interconnect_1:lpddr2_mp_cmd_reset_n_1_reset_bridge_in_reset_reset, mm_interconnect_1:video_dma_reset_n_reset_bridge_in_reset_reset, mm_interconnect_2:lpddr2_mp_cmd_reset_n_2_reset_bridge_in_reset_reset, mm_interconnect_2:mdma_from_idct_accel_reset_n_reset_bridge_in_reset_reset, mutex_0:reset_n, rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in0, rst_controller_003:reset_in0, sram:reset_reset, sram_bridge:reset, sram_sharer:reset_reset, sysid:reset_n, timer_0_0:reset_n, timer_0_1:reset_n, timer_1_0:reset_n, timer_1_1:reset_n, video_dma:reset_n_reset_n, video_fifo:wrreset_n, video_pll:rst, ycbcr_to_rgb_accelerator:reset_n]
	wire          sram_sharer_tcm_request;                                                      // sram_sharer:request -> sram_bridge:request
	wire    [1:0] sram_sharer_tcm_sram_tcm_byteenable_n_out_out;                                // sram_sharer:sram_tcm_byteenable_n_out -> sram_bridge:tcs_sram_tcm_byteenable_n_out
	wire          sram_sharer_tcm_sram_tcm_data_out_outen;                                      // sram_sharer:sram_tcm_data_outen -> sram_bridge:tcs_sram_tcm_data_outen
	wire   [15:0] sram_sharer_tcm_sram_tcm_data_out_in;                                         // sram_bridge:tcs_sram_tcm_data_in -> sram_sharer:sram_tcm_data_in
	wire    [0:0] sram_sharer_tcm_sram_tcm_write_n_out_out;                                     // sram_sharer:sram_tcm_write_n_out -> sram_bridge:tcs_sram_tcm_write_n_out
	wire   [15:0] sram_sharer_tcm_sram_tcm_data_out_out;                                        // sram_sharer:sram_tcm_data_out -> sram_bridge:tcs_sram_tcm_data_out
	wire   [18:0] sram_sharer_tcm_sram_tcm_address_out_out;                                     // sram_sharer:sram_tcm_address_out -> sram_bridge:tcs_sram_tcm_address_out
	wire    [0:0] sram_sharer_tcm_sram_tcm_chipselect_n_out_out;                                // sram_sharer:sram_tcm_chipselect_n_out -> sram_bridge:tcs_sram_tcm_chipselect_n_out
	wire          sram_sharer_tcm_grant;                                                        // sram_bridge:grant -> sram_sharer:grant
	wire    [0:0] sram_sharer_tcm_sram_tcm_outputenable_n_out_out;                              // sram_sharer:sram_tcm_outputenable_n_out -> sram_bridge:tcs_sram_tcm_outputenable_n_out
	wire          sram_tcm_data_outen;                                                          // sram:tcm_data_outen -> sram_sharer:tcs0_data_outen
	wire          sram_tcm_outputenable_n_out;                                                  // sram:tcm_outputenable_n_out -> sram_sharer:tcs0_outputenable_n_out
	wire          sram_tcm_request;                                                             // sram:tcm_request -> sram_sharer:tcs0_request
	wire    [1:0] sram_tcm_byteenable_n_out;                                                    // sram:tcm_byteenable_n_out -> sram_sharer:tcs0_byteenable_n_out
	wire          sram_tcm_write_n_out;                                                         // sram:tcm_write_n_out -> sram_sharer:tcs0_write_n_out
	wire          sram_tcm_grant;                                                               // sram_sharer:tcs0_grant -> sram:tcm_grant
	wire          sram_tcm_chipselect_n_out;                                                    // sram:tcm_chipselect_n_out -> sram_sharer:tcs0_chipselect_n_out
	wire   [18:0] sram_tcm_address_out;                                                         // sram:tcm_address_out -> sram_sharer:tcs0_address_out
	wire   [15:0] sram_tcm_data_out;                                                            // sram:tcm_data_out -> sram_sharer:tcs0_data_out
	wire   [15:0] sram_tcm_data_in;                                                             // sram_sharer:tcs0_data_in -> sram:tcm_data_in
	wire   [31:0] cpu_0_data_master_readdata;                                                   // mm_interconnect_0:cpu_0_data_master_readdata -> cpu_0:d_readdata
	wire          cpu_0_data_master_waitrequest;                                                // mm_interconnect_0:cpu_0_data_master_waitrequest -> cpu_0:d_waitrequest
	wire          cpu_0_data_master_debugaccess;                                                // cpu_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_0_data_master_debugaccess
	wire   [29:0] cpu_0_data_master_address;                                                    // cpu_0:d_address -> mm_interconnect_0:cpu_0_data_master_address
	wire    [3:0] cpu_0_data_master_byteenable;                                                 // cpu_0:d_byteenable -> mm_interconnect_0:cpu_0_data_master_byteenable
	wire          cpu_0_data_master_read;                                                       // cpu_0:d_read -> mm_interconnect_0:cpu_0_data_master_read
	wire          cpu_0_data_master_readdatavalid;                                              // mm_interconnect_0:cpu_0_data_master_readdatavalid -> cpu_0:d_readdatavalid
	wire          cpu_0_data_master_write;                                                      // cpu_0:d_write -> mm_interconnect_0:cpu_0_data_master_write
	wire   [31:0] cpu_0_data_master_writedata;                                                  // cpu_0:d_writedata -> mm_interconnect_0:cpu_0_data_master_writedata
	wire    [3:0] cpu_0_data_master_burstcount;                                                 // cpu_0:d_burstcount -> mm_interconnect_0:cpu_0_data_master_burstcount
	wire   [31:0] cpu_1_data_master_readdata;                                                   // mm_interconnect_0:cpu_1_data_master_readdata -> cpu_1:d_readdata
	wire          cpu_1_data_master_waitrequest;                                                // mm_interconnect_0:cpu_1_data_master_waitrequest -> cpu_1:d_waitrequest
	wire          cpu_1_data_master_debugaccess;                                                // cpu_1:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_1_data_master_debugaccess
	wire   [29:0] cpu_1_data_master_address;                                                    // cpu_1:d_address -> mm_interconnect_0:cpu_1_data_master_address
	wire    [3:0] cpu_1_data_master_byteenable;                                                 // cpu_1:d_byteenable -> mm_interconnect_0:cpu_1_data_master_byteenable
	wire          cpu_1_data_master_read;                                                       // cpu_1:d_read -> mm_interconnect_0:cpu_1_data_master_read
	wire          cpu_1_data_master_readdatavalid;                                              // mm_interconnect_0:cpu_1_data_master_readdatavalid -> cpu_1:d_readdatavalid
	wire          cpu_1_data_master_write;                                                      // cpu_1:d_write -> mm_interconnect_0:cpu_1_data_master_write
	wire   [31:0] cpu_1_data_master_writedata;                                                  // cpu_1:d_writedata -> mm_interconnect_0:cpu_1_data_master_writedata
	wire    [3:0] cpu_1_data_master_burstcount;                                                 // cpu_1:d_burstcount -> mm_interconnect_0:cpu_1_data_master_burstcount
	wire   [31:0] cpu_0_instruction_master_readdata;                                            // mm_interconnect_0:cpu_0_instruction_master_readdata -> cpu_0:i_readdata
	wire          cpu_0_instruction_master_waitrequest;                                         // mm_interconnect_0:cpu_0_instruction_master_waitrequest -> cpu_0:i_waitrequest
	wire   [29:0] cpu_0_instruction_master_address;                                             // cpu_0:i_address -> mm_interconnect_0:cpu_0_instruction_master_address
	wire          cpu_0_instruction_master_read;                                                // cpu_0:i_read -> mm_interconnect_0:cpu_0_instruction_master_read
	wire          cpu_0_instruction_master_readdatavalid;                                       // mm_interconnect_0:cpu_0_instruction_master_readdatavalid -> cpu_0:i_readdatavalid
	wire   [31:0] cpu_1_instruction_master_readdata;                                            // mm_interconnect_0:cpu_1_instruction_master_readdata -> cpu_1:i_readdata
	wire          cpu_1_instruction_master_waitrequest;                                         // mm_interconnect_0:cpu_1_instruction_master_waitrequest -> cpu_1:i_waitrequest
	wire   [29:0] cpu_1_instruction_master_address;                                             // cpu_1:i_address -> mm_interconnect_0:cpu_1_instruction_master_address
	wire          cpu_1_instruction_master_read;                                                // cpu_1:i_read -> mm_interconnect_0:cpu_1_instruction_master_read
	wire          cpu_1_instruction_master_readdatavalid;                                       // mm_interconnect_0:cpu_1_instruction_master_readdatavalid -> cpu_1:i_readdatavalid
	wire   [31:0] sd_cont_master_readdata;                                                      // mm_interconnect_0:sd_cont_master_readdata -> sd_cont:m_readdata
	wire          sd_cont_master_waitrequest;                                                   // mm_interconnect_0:sd_cont_master_waitrequest -> sd_cont:m_waitrequest_n
	wire   [31:0] sd_cont_master_address;                                                       // sd_cont:m_address -> mm_interconnect_0:sd_cont_master_address
	wire          sd_cont_master_read;                                                          // sd_cont:m_read -> mm_interconnect_0:sd_cont_master_read
	wire          sd_cont_master_write;                                                         // sd_cont:m_write -> mm_interconnect_0:sd_cont_master_write
	wire   [31:0] sd_cont_master_writedata;                                                     // sd_cont:m_writedata -> mm_interconnect_0:sd_cont_master_writedata
	wire          mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;                   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire   [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;                     // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire          mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;                  // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire    [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;                      // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire          mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;                         // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire          mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;                        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire   [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;                    // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire          mm_interconnect_0_lpddr2_avl_0_beginbursttransfer;                            // mm_interconnect_0:lpddr2_avl_0_beginbursttransfer -> lpddr2:avl_burstbegin_0
	wire   [31:0] mm_interconnect_0_lpddr2_avl_0_readdata;                                      // lpddr2:avl_rdata_0 -> mm_interconnect_0:lpddr2_avl_0_readdata
	wire          mm_interconnect_0_lpddr2_avl_0_waitrequest;                                   // lpddr2:avl_ready_0 -> mm_interconnect_0:lpddr2_avl_0_waitrequest
	wire   [26:0] mm_interconnect_0_lpddr2_avl_0_address;                                       // mm_interconnect_0:lpddr2_avl_0_address -> lpddr2:avl_addr_0
	wire          mm_interconnect_0_lpddr2_avl_0_read;                                          // mm_interconnect_0:lpddr2_avl_0_read -> lpddr2:avl_read_req_0
	wire    [3:0] mm_interconnect_0_lpddr2_avl_0_byteenable;                                    // mm_interconnect_0:lpddr2_avl_0_byteenable -> lpddr2:avl_be_0
	wire          mm_interconnect_0_lpddr2_avl_0_readdatavalid;                                 // lpddr2:avl_rdata_valid_0 -> mm_interconnect_0:lpddr2_avl_0_readdatavalid
	wire          mm_interconnect_0_lpddr2_avl_0_write;                                         // mm_interconnect_0:lpddr2_avl_0_write -> lpddr2:avl_write_req_0
	wire   [31:0] mm_interconnect_0_lpddr2_avl_0_writedata;                                     // mm_interconnect_0:lpddr2_avl_0_writedata -> lpddr2:avl_wdata_0
	wire    [7:0] mm_interconnect_0_lpddr2_avl_0_burstcount;                                    // mm_interconnect_0:lpddr2_avl_0_burstcount -> lpddr2:avl_size_0
	wire   [31:0] mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_receiver_readdata;     // mailbox_simple_cpu1_to_cpu0:avmm_rcv_readdata -> mm_interconnect_0:mailbox_simple_cpu1_to_cpu0_avmm_msg_receiver_readdata
	wire    [1:0] mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_receiver_address;      // mm_interconnect_0:mailbox_simple_cpu1_to_cpu0_avmm_msg_receiver_address -> mailbox_simple_cpu1_to_cpu0:avmm_rcv_address
	wire          mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_receiver_read;         // mm_interconnect_0:mailbox_simple_cpu1_to_cpu0_avmm_msg_receiver_read -> mailbox_simple_cpu1_to_cpu0:avmm_rcv_read
	wire          mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_receiver_write;        // mm_interconnect_0:mailbox_simple_cpu1_to_cpu0_avmm_msg_receiver_write -> mailbox_simple_cpu1_to_cpu0:avmm_rcv_write
	wire   [31:0] mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_receiver_writedata;    // mm_interconnect_0:mailbox_simple_cpu1_to_cpu0_avmm_msg_receiver_writedata -> mailbox_simple_cpu1_to_cpu0:avmm_rcv_writedata
	wire   [31:0] mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_sender_readdata;       // mailbox_simple_cpu0_to_cpu1:avmm_snd_readdata -> mm_interconnect_0:mailbox_simple_cpu0_to_cpu1_avmm_msg_sender_readdata
	wire          mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_sender_waitrequest;    // mailbox_simple_cpu0_to_cpu1:avmm_snd_waitrequest -> mm_interconnect_0:mailbox_simple_cpu0_to_cpu1_avmm_msg_sender_waitrequest
	wire    [1:0] mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_sender_address;        // mm_interconnect_0:mailbox_simple_cpu0_to_cpu1_avmm_msg_sender_address -> mailbox_simple_cpu0_to_cpu1:avmm_snd_address
	wire          mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_sender_read;           // mm_interconnect_0:mailbox_simple_cpu0_to_cpu1_avmm_msg_sender_read -> mailbox_simple_cpu0_to_cpu1:avmm_snd_read
	wire          mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_sender_write;          // mm_interconnect_0:mailbox_simple_cpu0_to_cpu1_avmm_msg_sender_write -> mailbox_simple_cpu0_to_cpu1:avmm_snd_write
	wire   [31:0] mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_sender_writedata;      // mm_interconnect_0:mailbox_simple_cpu0_to_cpu1_avmm_msg_sender_writedata -> mailbox_simple_cpu0_to_cpu1:avmm_snd_writedata
	wire   [31:0] mm_interconnect_0_sysid_control_slave_readdata;                               // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire    [0:0] mm_interconnect_0_sysid_control_slave_address;                                // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire   [31:0] mm_interconnect_0_video_dma_csr_readdata;                                     // video_dma:csr_readdata -> mm_interconnect_0:video_dma_csr_readdata
	wire    [2:0] mm_interconnect_0_video_dma_csr_address;                                      // mm_interconnect_0:video_dma_csr_address -> video_dma:csr_address
	wire          mm_interconnect_0_video_dma_csr_read;                                         // mm_interconnect_0:video_dma_csr_read -> video_dma:csr_read
	wire    [3:0] mm_interconnect_0_video_dma_csr_byteenable;                                   // mm_interconnect_0:video_dma_csr_byteenable -> video_dma:csr_byteenable
	wire          mm_interconnect_0_video_dma_csr_write;                                        // mm_interconnect_0:video_dma_csr_write -> video_dma:csr_write
	wire   [31:0] mm_interconnect_0_video_dma_csr_writedata;                                    // mm_interconnect_0:video_dma_csr_writedata -> video_dma:csr_writedata
	wire   [31:0] mm_interconnect_0_cpu_0_debug_mem_slave_readdata;                             // cpu_0:debug_mem_slave_readdata -> mm_interconnect_0:cpu_0_debug_mem_slave_readdata
	wire          mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest;                          // cpu_0:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_0_debug_mem_slave_waitrequest
	wire          mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess;                          // mm_interconnect_0:cpu_0_debug_mem_slave_debugaccess -> cpu_0:debug_mem_slave_debugaccess
	wire    [8:0] mm_interconnect_0_cpu_0_debug_mem_slave_address;                              // mm_interconnect_0:cpu_0_debug_mem_slave_address -> cpu_0:debug_mem_slave_address
	wire          mm_interconnect_0_cpu_0_debug_mem_slave_read;                                 // mm_interconnect_0:cpu_0_debug_mem_slave_read -> cpu_0:debug_mem_slave_read
	wire    [3:0] mm_interconnect_0_cpu_0_debug_mem_slave_byteenable;                           // mm_interconnect_0:cpu_0_debug_mem_slave_byteenable -> cpu_0:debug_mem_slave_byteenable
	wire          mm_interconnect_0_cpu_0_debug_mem_slave_write;                                // mm_interconnect_0:cpu_0_debug_mem_slave_write -> cpu_0:debug_mem_slave_write
	wire   [31:0] mm_interconnect_0_cpu_0_debug_mem_slave_writedata;                            // mm_interconnect_0:cpu_0_debug_mem_slave_writedata -> cpu_0:debug_mem_slave_writedata
	wire          mm_interconnect_0_video_dma_descriptor_slave_waitrequest;                     // video_dma:descriptor_slave_waitrequest -> mm_interconnect_0:video_dma_descriptor_slave_waitrequest
	wire   [15:0] mm_interconnect_0_video_dma_descriptor_slave_byteenable;                      // mm_interconnect_0:video_dma_descriptor_slave_byteenable -> video_dma:descriptor_slave_byteenable
	wire          mm_interconnect_0_video_dma_descriptor_slave_write;                           // mm_interconnect_0:video_dma_descriptor_slave_write -> video_dma:descriptor_slave_write
	wire  [127:0] mm_interconnect_0_video_dma_descriptor_slave_writedata;                       // mm_interconnect_0:video_dma_descriptor_slave_writedata -> video_dma:descriptor_slave_writedata
	wire          mm_interconnect_0_timer_0_0_s1_chipselect;                                    // mm_interconnect_0:timer_0_0_s1_chipselect -> timer_0_0:chipselect
	wire   [15:0] mm_interconnect_0_timer_0_0_s1_readdata;                                      // timer_0_0:readdata -> mm_interconnect_0:timer_0_0_s1_readdata
	wire    [2:0] mm_interconnect_0_timer_0_0_s1_address;                                       // mm_interconnect_0:timer_0_0_s1_address -> timer_0_0:address
	wire          mm_interconnect_0_timer_0_0_s1_write;                                         // mm_interconnect_0:timer_0_0_s1_write -> timer_0_0:write_n
	wire   [15:0] mm_interconnect_0_timer_0_0_s1_writedata;                                     // mm_interconnect_0:timer_0_0_s1_writedata -> timer_0_0:writedata
	wire          mm_interconnect_0_key_s1_chipselect;                                          // mm_interconnect_0:key_s1_chipselect -> key:chipselect
	wire   [31:0] mm_interconnect_0_key_s1_readdata;                                            // key:readdata -> mm_interconnect_0:key_s1_readdata
	wire    [1:0] mm_interconnect_0_key_s1_address;                                             // mm_interconnect_0:key_s1_address -> key:address
	wire          mm_interconnect_0_key_s1_write;                                               // mm_interconnect_0:key_s1_write -> key:write_n
	wire   [31:0] mm_interconnect_0_key_s1_writedata;                                           // mm_interconnect_0:key_s1_writedata -> key:writedata
	wire          mm_interconnect_0_timer_0_1_s1_chipselect;                                    // mm_interconnect_0:timer_0_1_s1_chipselect -> timer_0_1:chipselect
	wire   [15:0] mm_interconnect_0_timer_0_1_s1_readdata;                                      // timer_0_1:readdata -> mm_interconnect_0:timer_0_1_s1_readdata
	wire    [3:0] mm_interconnect_0_timer_0_1_s1_address;                                       // mm_interconnect_0:timer_0_1_s1_address -> timer_0_1:address
	wire          mm_interconnect_0_timer_0_1_s1_write;                                         // mm_interconnect_0:timer_0_1_s1_write -> timer_0_1:write_n
	wire   [15:0] mm_interconnect_0_timer_0_1_s1_writedata;                                     // mm_interconnect_0:timer_0_1_s1_writedata -> timer_0_1:writedata
	wire          mm_interconnect_0_ledg_s1_chipselect;                                         // mm_interconnect_0:ledg_s1_chipselect -> ledg:chipselect
	wire   [31:0] mm_interconnect_0_ledg_s1_readdata;                                           // ledg:readdata -> mm_interconnect_0:ledg_s1_readdata
	wire    [2:0] mm_interconnect_0_ledg_s1_address;                                            // mm_interconnect_0:ledg_s1_address -> ledg:address
	wire          mm_interconnect_0_ledg_s1_write;                                              // mm_interconnect_0:ledg_s1_write -> ledg:write_n
	wire   [31:0] mm_interconnect_0_ledg_s1_writedata;                                          // mm_interconnect_0:ledg_s1_writedata -> ledg:writedata
	wire          mm_interconnect_0_ledr_s1_chipselect;                                         // mm_interconnect_0:ledr_s1_chipselect -> ledr:chipselect
	wire   [31:0] mm_interconnect_0_ledr_s1_readdata;                                           // ledr:readdata -> mm_interconnect_0:ledr_s1_readdata
	wire    [2:0] mm_interconnect_0_ledr_s1_address;                                            // mm_interconnect_0:ledr_s1_address -> ledr:address
	wire          mm_interconnect_0_ledr_s1_write;                                              // mm_interconnect_0:ledr_s1_write -> ledr:write_n
	wire   [31:0] mm_interconnect_0_ledr_s1_writedata;                                          // mm_interconnect_0:ledr_s1_writedata -> ledr:writedata
	wire          mm_interconnect_0_i2c_scl_s1_chipselect;                                      // mm_interconnect_0:i2c_scl_s1_chipselect -> i2c_scl:chipselect
	wire   [31:0] mm_interconnect_0_i2c_scl_s1_readdata;                                        // i2c_scl:readdata -> mm_interconnect_0:i2c_scl_s1_readdata
	wire    [1:0] mm_interconnect_0_i2c_scl_s1_address;                                         // mm_interconnect_0:i2c_scl_s1_address -> i2c_scl:address
	wire          mm_interconnect_0_i2c_scl_s1_write;                                           // mm_interconnect_0:i2c_scl_s1_write -> i2c_scl:write_n
	wire   [31:0] mm_interconnect_0_i2c_scl_s1_writedata;                                       // mm_interconnect_0:i2c_scl_s1_writedata -> i2c_scl:writedata
	wire          mm_interconnect_0_i2c_sda_s1_chipselect;                                      // mm_interconnect_0:i2c_sda_s1_chipselect -> i2c_sda:chipselect
	wire   [31:0] mm_interconnect_0_i2c_sda_s1_readdata;                                        // i2c_sda:readdata -> mm_interconnect_0:i2c_sda_s1_readdata
	wire    [1:0] mm_interconnect_0_i2c_sda_s1_address;                                         // mm_interconnect_0:i2c_sda_s1_address -> i2c_sda:address
	wire          mm_interconnect_0_i2c_sda_s1_write;                                           // mm_interconnect_0:i2c_sda_s1_write -> i2c_sda:write_n
	wire   [31:0] mm_interconnect_0_i2c_sda_s1_writedata;                                       // mm_interconnect_0:i2c_sda_s1_writedata -> i2c_sda:writedata
	wire          mm_interconnect_0_mutex_0_s1_chipselect;                                      // mm_interconnect_0:mutex_0_s1_chipselect -> mutex_0:chipselect
	wire   [31:0] mm_interconnect_0_mutex_0_s1_readdata;                                        // mutex_0:data_to_cpu -> mm_interconnect_0:mutex_0_s1_readdata
	wire    [0:0] mm_interconnect_0_mutex_0_s1_address;                                         // mm_interconnect_0:mutex_0_s1_address -> mutex_0:address
	wire          mm_interconnect_0_mutex_0_s1_read;                                            // mm_interconnect_0:mutex_0_s1_read -> mutex_0:read
	wire          mm_interconnect_0_mutex_0_s1_write;                                           // mm_interconnect_0:mutex_0_s1_write -> mutex_0:write
	wire   [31:0] mm_interconnect_0_mutex_0_s1_writedata;                                       // mm_interconnect_0:mutex_0_s1_writedata -> mutex_0:data_from_cpu
	wire          mm_interconnect_0_sd_cont_slave_chipselect;                                   // mm_interconnect_0:sd_cont_slave_chipselect -> sd_cont:s_chipselect
	wire   [31:0] mm_interconnect_0_sd_cont_slave_readdata;                                     // sd_cont:s_readdata -> mm_interconnect_0:sd_cont_slave_readdata
	wire          mm_interconnect_0_sd_cont_slave_waitrequest;                                  // sd_cont:s_waitrequest_n -> mm_interconnect_0:sd_cont_slave_waitrequest
	wire    [7:0] mm_interconnect_0_sd_cont_slave_address;                                      // mm_interconnect_0:sd_cont_slave_address -> sd_cont:s_address
	wire          mm_interconnect_0_sd_cont_slave_read;                                         // mm_interconnect_0:sd_cont_slave_read -> sd_cont:s_read
	wire          mm_interconnect_0_sd_cont_slave_write;                                        // mm_interconnect_0:sd_cont_slave_write -> sd_cont:s_write
	wire   [31:0] mm_interconnect_0_sd_cont_slave_writedata;                                    // mm_interconnect_0:sd_cont_slave_writedata -> sd_cont:s_writedata
	wire   [15:0] mm_interconnect_0_sram_uas_readdata;                                          // sram:uas_readdata -> mm_interconnect_0:sram_uas_readdata
	wire          mm_interconnect_0_sram_uas_waitrequest;                                       // sram:uas_waitrequest -> mm_interconnect_0:sram_uas_waitrequest
	wire          mm_interconnect_0_sram_uas_debugaccess;                                       // mm_interconnect_0:sram_uas_debugaccess -> sram:uas_debugaccess
	wire   [18:0] mm_interconnect_0_sram_uas_address;                                           // mm_interconnect_0:sram_uas_address -> sram:uas_address
	wire          mm_interconnect_0_sram_uas_read;                                              // mm_interconnect_0:sram_uas_read -> sram:uas_read
	wire    [1:0] mm_interconnect_0_sram_uas_byteenable;                                        // mm_interconnect_0:sram_uas_byteenable -> sram:uas_byteenable
	wire          mm_interconnect_0_sram_uas_readdatavalid;                                     // sram:uas_readdatavalid -> mm_interconnect_0:sram_uas_readdatavalid
	wire          mm_interconnect_0_sram_uas_lock;                                              // mm_interconnect_0:sram_uas_lock -> sram:uas_lock
	wire          mm_interconnect_0_sram_uas_write;                                             // mm_interconnect_0:sram_uas_write -> sram:uas_write
	wire   [15:0] mm_interconnect_0_sram_uas_writedata;                                         // mm_interconnect_0:sram_uas_writedata -> sram:uas_writedata
	wire    [1:0] mm_interconnect_0_sram_uas_burstcount;                                        // mm_interconnect_0:sram_uas_burstcount -> sram:uas_burstcount
	wire   [31:0] mm_interconnect_0_cpu_1_debug_mem_slave_readdata;                             // cpu_1:debug_mem_slave_readdata -> mm_interconnect_0:cpu_1_debug_mem_slave_readdata
	wire          mm_interconnect_0_cpu_1_debug_mem_slave_waitrequest;                          // cpu_1:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_1_debug_mem_slave_waitrequest
	wire          mm_interconnect_0_cpu_1_debug_mem_slave_debugaccess;                          // mm_interconnect_0:cpu_1_debug_mem_slave_debugaccess -> cpu_1:debug_mem_slave_debugaccess
	wire    [8:0] mm_interconnect_0_cpu_1_debug_mem_slave_address;                              // mm_interconnect_0:cpu_1_debug_mem_slave_address -> cpu_1:debug_mem_slave_address
	wire          mm_interconnect_0_cpu_1_debug_mem_slave_read;                                 // mm_interconnect_0:cpu_1_debug_mem_slave_read -> cpu_1:debug_mem_slave_read
	wire    [3:0] mm_interconnect_0_cpu_1_debug_mem_slave_byteenable;                           // mm_interconnect_0:cpu_1_debug_mem_slave_byteenable -> cpu_1:debug_mem_slave_byteenable
	wire          mm_interconnect_0_cpu_1_debug_mem_slave_write;                                // mm_interconnect_0:cpu_1_debug_mem_slave_write -> cpu_1:debug_mem_slave_write
	wire   [31:0] mm_interconnect_0_cpu_1_debug_mem_slave_writedata;                            // mm_interconnect_0:cpu_1_debug_mem_slave_writedata -> cpu_1:debug_mem_slave_writedata
	wire          mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_chipselect;                   // mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_chipselect -> jtag_uart_1:av_chipselect
	wire   [31:0] mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_readdata;                     // jtag_uart_1:av_readdata -> mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_readdata
	wire          mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_waitrequest;                  // jtag_uart_1:av_waitrequest -> mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_waitrequest
	wire    [0:0] mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_address;                      // mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_address -> jtag_uart_1:av_address
	wire          mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read;                         // mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_read -> jtag_uart_1:av_read_n
	wire          mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write;                        // mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_write -> jtag_uart_1:av_write_n
	wire   [31:0] mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_writedata;                    // mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_writedata -> jtag_uart_1:av_writedata
	wire   [31:0] mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_receiver_readdata;     // mailbox_simple_cpu0_to_cpu1:avmm_rcv_readdata -> mm_interconnect_0:mailbox_simple_cpu0_to_cpu1_avmm_msg_receiver_readdata
	wire    [1:0] mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_receiver_address;      // mm_interconnect_0:mailbox_simple_cpu0_to_cpu1_avmm_msg_receiver_address -> mailbox_simple_cpu0_to_cpu1:avmm_rcv_address
	wire          mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_receiver_read;         // mm_interconnect_0:mailbox_simple_cpu0_to_cpu1_avmm_msg_receiver_read -> mailbox_simple_cpu0_to_cpu1:avmm_rcv_read
	wire          mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_receiver_write;        // mm_interconnect_0:mailbox_simple_cpu0_to_cpu1_avmm_msg_receiver_write -> mailbox_simple_cpu0_to_cpu1:avmm_rcv_write
	wire   [31:0] mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_receiver_writedata;    // mm_interconnect_0:mailbox_simple_cpu0_to_cpu1_avmm_msg_receiver_writedata -> mailbox_simple_cpu0_to_cpu1:avmm_rcv_writedata
	wire   [31:0] mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_sender_readdata;       // mailbox_simple_cpu1_to_cpu0:avmm_snd_readdata -> mm_interconnect_0:mailbox_simple_cpu1_to_cpu0_avmm_msg_sender_readdata
	wire          mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_sender_waitrequest;    // mailbox_simple_cpu1_to_cpu0:avmm_snd_waitrequest -> mm_interconnect_0:mailbox_simple_cpu1_to_cpu0_avmm_msg_sender_waitrequest
	wire    [1:0] mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_sender_address;        // mm_interconnect_0:mailbox_simple_cpu1_to_cpu0_avmm_msg_sender_address -> mailbox_simple_cpu1_to_cpu0:avmm_snd_address
	wire          mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_sender_read;           // mm_interconnect_0:mailbox_simple_cpu1_to_cpu0_avmm_msg_sender_read -> mailbox_simple_cpu1_to_cpu0:avmm_snd_read
	wire          mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_sender_write;          // mm_interconnect_0:mailbox_simple_cpu1_to_cpu0_avmm_msg_sender_write -> mailbox_simple_cpu1_to_cpu0:avmm_snd_write
	wire   [31:0] mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_sender_writedata;      // mm_interconnect_0:mailbox_simple_cpu1_to_cpu0_avmm_msg_sender_writedata -> mailbox_simple_cpu1_to_cpu0:avmm_snd_writedata
	wire   [31:0] mm_interconnect_0_mdma_to_idct_accel_csr_readdata;                            // mdma_to_idct_accel:csr_readdata -> mm_interconnect_0:mdma_to_idct_accel_csr_readdata
	wire    [2:0] mm_interconnect_0_mdma_to_idct_accel_csr_address;                             // mm_interconnect_0:mdma_to_idct_accel_csr_address -> mdma_to_idct_accel:csr_address
	wire          mm_interconnect_0_mdma_to_idct_accel_csr_read;                                // mm_interconnect_0:mdma_to_idct_accel_csr_read -> mdma_to_idct_accel:csr_read
	wire    [3:0] mm_interconnect_0_mdma_to_idct_accel_csr_byteenable;                          // mm_interconnect_0:mdma_to_idct_accel_csr_byteenable -> mdma_to_idct_accel:csr_byteenable
	wire          mm_interconnect_0_mdma_to_idct_accel_csr_write;                               // mm_interconnect_0:mdma_to_idct_accel_csr_write -> mdma_to_idct_accel:csr_write
	wire   [31:0] mm_interconnect_0_mdma_to_idct_accel_csr_writedata;                           // mm_interconnect_0:mdma_to_idct_accel_csr_writedata -> mdma_to_idct_accel:csr_writedata
	wire   [31:0] mm_interconnect_0_mdma_from_idct_accel_csr_readdata;                          // mdma_from_idct_accel:csr_readdata -> mm_interconnect_0:mdma_from_idct_accel_csr_readdata
	wire    [2:0] mm_interconnect_0_mdma_from_idct_accel_csr_address;                           // mm_interconnect_0:mdma_from_idct_accel_csr_address -> mdma_from_idct_accel:csr_address
	wire          mm_interconnect_0_mdma_from_idct_accel_csr_read;                              // mm_interconnect_0:mdma_from_idct_accel_csr_read -> mdma_from_idct_accel:csr_read
	wire    [3:0] mm_interconnect_0_mdma_from_idct_accel_csr_byteenable;                        // mm_interconnect_0:mdma_from_idct_accel_csr_byteenable -> mdma_from_idct_accel:csr_byteenable
	wire          mm_interconnect_0_mdma_from_idct_accel_csr_write;                             // mm_interconnect_0:mdma_from_idct_accel_csr_write -> mdma_from_idct_accel:csr_write
	wire   [31:0] mm_interconnect_0_mdma_from_idct_accel_csr_writedata;                         // mm_interconnect_0:mdma_from_idct_accel_csr_writedata -> mdma_from_idct_accel:csr_writedata
	wire   [31:0] mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cb_csr_readdata;                 // mdma_to_ycbcr_to_rgb_accel_cb:csr_readdata -> mm_interconnect_0:mdma_to_ycbcr_to_rgb_accel_cb_csr_readdata
	wire    [2:0] mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cb_csr_address;                  // mm_interconnect_0:mdma_to_ycbcr_to_rgb_accel_cb_csr_address -> mdma_to_ycbcr_to_rgb_accel_cb:csr_address
	wire          mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cb_csr_read;                     // mm_interconnect_0:mdma_to_ycbcr_to_rgb_accel_cb_csr_read -> mdma_to_ycbcr_to_rgb_accel_cb:csr_read
	wire    [3:0] mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cb_csr_byteenable;               // mm_interconnect_0:mdma_to_ycbcr_to_rgb_accel_cb_csr_byteenable -> mdma_to_ycbcr_to_rgb_accel_cb:csr_byteenable
	wire          mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cb_csr_write;                    // mm_interconnect_0:mdma_to_ycbcr_to_rgb_accel_cb_csr_write -> mdma_to_ycbcr_to_rgb_accel_cb:csr_write
	wire   [31:0] mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cb_csr_writedata;                // mm_interconnect_0:mdma_to_ycbcr_to_rgb_accel_cb_csr_writedata -> mdma_to_ycbcr_to_rgb_accel_cb:csr_writedata
	wire   [31:0] mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cr_csr_readdata;                 // mdma_to_ycbcr_to_rgb_accel_cr:csr_readdata -> mm_interconnect_0:mdma_to_ycbcr_to_rgb_accel_cr_csr_readdata
	wire    [2:0] mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cr_csr_address;                  // mm_interconnect_0:mdma_to_ycbcr_to_rgb_accel_cr_csr_address -> mdma_to_ycbcr_to_rgb_accel_cr:csr_address
	wire          mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cr_csr_read;                     // mm_interconnect_0:mdma_to_ycbcr_to_rgb_accel_cr_csr_read -> mdma_to_ycbcr_to_rgb_accel_cr:csr_read
	wire    [3:0] mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cr_csr_byteenable;               // mm_interconnect_0:mdma_to_ycbcr_to_rgb_accel_cr_csr_byteenable -> mdma_to_ycbcr_to_rgb_accel_cr:csr_byteenable
	wire          mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cr_csr_write;                    // mm_interconnect_0:mdma_to_ycbcr_to_rgb_accel_cr_csr_write -> mdma_to_ycbcr_to_rgb_accel_cr:csr_write
	wire   [31:0] mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cr_csr_writedata;                // mm_interconnect_0:mdma_to_ycbcr_to_rgb_accel_cr_csr_writedata -> mdma_to_ycbcr_to_rgb_accel_cr:csr_writedata
	wire   [31:0] mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_y_csr_readdata;                  // mdma_to_ycbcr_to_rgb_accel_y:csr_readdata -> mm_interconnect_0:mdma_to_ycbcr_to_rgb_accel_y_csr_readdata
	wire    [2:0] mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_y_csr_address;                   // mm_interconnect_0:mdma_to_ycbcr_to_rgb_accel_y_csr_address -> mdma_to_ycbcr_to_rgb_accel_y:csr_address
	wire          mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_y_csr_read;                      // mm_interconnect_0:mdma_to_ycbcr_to_rgb_accel_y_csr_read -> mdma_to_ycbcr_to_rgb_accel_y:csr_read
	wire    [3:0] mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_y_csr_byteenable;                // mm_interconnect_0:mdma_to_ycbcr_to_rgb_accel_y_csr_byteenable -> mdma_to_ycbcr_to_rgb_accel_y:csr_byteenable
	wire          mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_y_csr_write;                     // mm_interconnect_0:mdma_to_ycbcr_to_rgb_accel_y_csr_write -> mdma_to_ycbcr_to_rgb_accel_y:csr_write
	wire   [31:0] mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_y_csr_writedata;                 // mm_interconnect_0:mdma_to_ycbcr_to_rgb_accel_y_csr_writedata -> mdma_to_ycbcr_to_rgb_accel_y:csr_writedata
	wire   [31:0] mm_interconnect_0_mdma_from_ycbcr_to_rgb_accel_csr_readdata;                  // mdma_from_ycbcr_to_rgb_accel:csr_readdata -> mm_interconnect_0:mdma_from_ycbcr_to_rgb_accel_csr_readdata
	wire    [2:0] mm_interconnect_0_mdma_from_ycbcr_to_rgb_accel_csr_address;                   // mm_interconnect_0:mdma_from_ycbcr_to_rgb_accel_csr_address -> mdma_from_ycbcr_to_rgb_accel:csr_address
	wire          mm_interconnect_0_mdma_from_ycbcr_to_rgb_accel_csr_read;                      // mm_interconnect_0:mdma_from_ycbcr_to_rgb_accel_csr_read -> mdma_from_ycbcr_to_rgb_accel:csr_read
	wire    [3:0] mm_interconnect_0_mdma_from_ycbcr_to_rgb_accel_csr_byteenable;                // mm_interconnect_0:mdma_from_ycbcr_to_rgb_accel_csr_byteenable -> mdma_from_ycbcr_to_rgb_accel:csr_byteenable
	wire          mm_interconnect_0_mdma_from_ycbcr_to_rgb_accel_csr_write;                     // mm_interconnect_0:mdma_from_ycbcr_to_rgb_accel_csr_write -> mdma_from_ycbcr_to_rgb_accel:csr_write
	wire   [31:0] mm_interconnect_0_mdma_from_ycbcr_to_rgb_accel_csr_writedata;                 // mm_interconnect_0:mdma_from_ycbcr_to_rgb_accel_csr_writedata -> mdma_from_ycbcr_to_rgb_accel:csr_writedata
	wire          mm_interconnect_0_mdma_to_idct_accel_descriptor_slave_waitrequest;            // mdma_to_idct_accel:descriptor_slave_waitrequest -> mm_interconnect_0:mdma_to_idct_accel_descriptor_slave_waitrequest
	wire   [15:0] mm_interconnect_0_mdma_to_idct_accel_descriptor_slave_byteenable;             // mm_interconnect_0:mdma_to_idct_accel_descriptor_slave_byteenable -> mdma_to_idct_accel:descriptor_slave_byteenable
	wire          mm_interconnect_0_mdma_to_idct_accel_descriptor_slave_write;                  // mm_interconnect_0:mdma_to_idct_accel_descriptor_slave_write -> mdma_to_idct_accel:descriptor_slave_write
	wire  [127:0] mm_interconnect_0_mdma_to_idct_accel_descriptor_slave_writedata;              // mm_interconnect_0:mdma_to_idct_accel_descriptor_slave_writedata -> mdma_to_idct_accel:descriptor_slave_writedata
	wire          mm_interconnect_0_mdma_from_idct_accel_descriptor_slave_waitrequest;          // mdma_from_idct_accel:descriptor_slave_waitrequest -> mm_interconnect_0:mdma_from_idct_accel_descriptor_slave_waitrequest
	wire   [15:0] mm_interconnect_0_mdma_from_idct_accel_descriptor_slave_byteenable;           // mm_interconnect_0:mdma_from_idct_accel_descriptor_slave_byteenable -> mdma_from_idct_accel:descriptor_slave_byteenable
	wire          mm_interconnect_0_mdma_from_idct_accel_descriptor_slave_write;                // mm_interconnect_0:mdma_from_idct_accel_descriptor_slave_write -> mdma_from_idct_accel:descriptor_slave_write
	wire  [127:0] mm_interconnect_0_mdma_from_idct_accel_descriptor_slave_writedata;            // mm_interconnect_0:mdma_from_idct_accel_descriptor_slave_writedata -> mdma_from_idct_accel:descriptor_slave_writedata
	wire          mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cb_descriptor_slave_waitrequest; // mdma_to_ycbcr_to_rgb_accel_cb:descriptor_slave_waitrequest -> mm_interconnect_0:mdma_to_ycbcr_to_rgb_accel_cb_descriptor_slave_waitrequest
	wire   [15:0] mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cb_descriptor_slave_byteenable;  // mm_interconnect_0:mdma_to_ycbcr_to_rgb_accel_cb_descriptor_slave_byteenable -> mdma_to_ycbcr_to_rgb_accel_cb:descriptor_slave_byteenable
	wire          mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cb_descriptor_slave_write;       // mm_interconnect_0:mdma_to_ycbcr_to_rgb_accel_cb_descriptor_slave_write -> mdma_to_ycbcr_to_rgb_accel_cb:descriptor_slave_write
	wire  [127:0] mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cb_descriptor_slave_writedata;   // mm_interconnect_0:mdma_to_ycbcr_to_rgb_accel_cb_descriptor_slave_writedata -> mdma_to_ycbcr_to_rgb_accel_cb:descriptor_slave_writedata
	wire          mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cr_descriptor_slave_waitrequest; // mdma_to_ycbcr_to_rgb_accel_cr:descriptor_slave_waitrequest -> mm_interconnect_0:mdma_to_ycbcr_to_rgb_accel_cr_descriptor_slave_waitrequest
	wire   [15:0] mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cr_descriptor_slave_byteenable;  // mm_interconnect_0:mdma_to_ycbcr_to_rgb_accel_cr_descriptor_slave_byteenable -> mdma_to_ycbcr_to_rgb_accel_cr:descriptor_slave_byteenable
	wire          mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cr_descriptor_slave_write;       // mm_interconnect_0:mdma_to_ycbcr_to_rgb_accel_cr_descriptor_slave_write -> mdma_to_ycbcr_to_rgb_accel_cr:descriptor_slave_write
	wire  [127:0] mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cr_descriptor_slave_writedata;   // mm_interconnect_0:mdma_to_ycbcr_to_rgb_accel_cr_descriptor_slave_writedata -> mdma_to_ycbcr_to_rgb_accel_cr:descriptor_slave_writedata
	wire          mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_y_descriptor_slave_waitrequest;  // mdma_to_ycbcr_to_rgb_accel_y:descriptor_slave_waitrequest -> mm_interconnect_0:mdma_to_ycbcr_to_rgb_accel_y_descriptor_slave_waitrequest
	wire   [15:0] mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_y_descriptor_slave_byteenable;   // mm_interconnect_0:mdma_to_ycbcr_to_rgb_accel_y_descriptor_slave_byteenable -> mdma_to_ycbcr_to_rgb_accel_y:descriptor_slave_byteenable
	wire          mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_y_descriptor_slave_write;        // mm_interconnect_0:mdma_to_ycbcr_to_rgb_accel_y_descriptor_slave_write -> mdma_to_ycbcr_to_rgb_accel_y:descriptor_slave_write
	wire  [127:0] mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_y_descriptor_slave_writedata;    // mm_interconnect_0:mdma_to_ycbcr_to_rgb_accel_y_descriptor_slave_writedata -> mdma_to_ycbcr_to_rgb_accel_y:descriptor_slave_writedata
	wire          mm_interconnect_0_mdma_from_ycbcr_to_rgb_accel_descriptor_slave_waitrequest;  // mdma_from_ycbcr_to_rgb_accel:descriptor_slave_waitrequest -> mm_interconnect_0:mdma_from_ycbcr_to_rgb_accel_descriptor_slave_waitrequest
	wire   [15:0] mm_interconnect_0_mdma_from_ycbcr_to_rgb_accel_descriptor_slave_byteenable;   // mm_interconnect_0:mdma_from_ycbcr_to_rgb_accel_descriptor_slave_byteenable -> mdma_from_ycbcr_to_rgb_accel:descriptor_slave_byteenable
	wire          mm_interconnect_0_mdma_from_ycbcr_to_rgb_accel_descriptor_slave_write;        // mm_interconnect_0:mdma_from_ycbcr_to_rgb_accel_descriptor_slave_write -> mdma_from_ycbcr_to_rgb_accel:descriptor_slave_write
	wire  [127:0] mm_interconnect_0_mdma_from_ycbcr_to_rgb_accel_descriptor_slave_writedata;    // mm_interconnect_0:mdma_from_ycbcr_to_rgb_accel_descriptor_slave_writedata -> mdma_from_ycbcr_to_rgb_accel:descriptor_slave_writedata
	wire          mm_interconnect_0_timer_1_0_s1_chipselect;                                    // mm_interconnect_0:timer_1_0_s1_chipselect -> timer_1_0:chipselect
	wire   [15:0] mm_interconnect_0_timer_1_0_s1_readdata;                                      // timer_1_0:readdata -> mm_interconnect_0:timer_1_0_s1_readdata
	wire    [3:0] mm_interconnect_0_timer_1_0_s1_address;                                       // mm_interconnect_0:timer_1_0_s1_address -> timer_1_0:address
	wire          mm_interconnect_0_timer_1_0_s1_write;                                         // mm_interconnect_0:timer_1_0_s1_write -> timer_1_0:write_n
	wire   [15:0] mm_interconnect_0_timer_1_0_s1_writedata;                                     // mm_interconnect_0:timer_1_0_s1_writedata -> timer_1_0:writedata
	wire          mm_interconnect_0_timer_1_1_s1_chipselect;                                    // mm_interconnect_0:timer_1_1_s1_chipselect -> timer_1_1:chipselect
	wire   [15:0] mm_interconnect_0_timer_1_1_s1_readdata;                                      // timer_1_1:readdata -> mm_interconnect_0:timer_1_1_s1_readdata
	wire    [3:0] mm_interconnect_0_timer_1_1_s1_address;                                       // mm_interconnect_0:timer_1_1_s1_address -> timer_1_1:address
	wire          mm_interconnect_0_timer_1_1_s1_write;                                         // mm_interconnect_0:timer_1_1_s1_write -> timer_1_1:write_n
	wire   [15:0] mm_interconnect_0_timer_1_1_s1_writedata;                                     // mm_interconnect_0:timer_1_1_s1_writedata -> timer_1_1:writedata
	wire   [31:0] video_dma_mm_read_readdata;                                                   // mm_interconnect_1:video_dma_mm_read_readdata -> video_dma:mm_read_readdata
	wire          video_dma_mm_read_waitrequest;                                                // mm_interconnect_1:video_dma_mm_read_waitrequest -> video_dma:mm_read_waitrequest
	wire   [28:0] video_dma_mm_read_address;                                                    // video_dma:mm_read_address -> mm_interconnect_1:video_dma_mm_read_address
	wire          video_dma_mm_read_read;                                                       // video_dma:mm_read_read -> mm_interconnect_1:video_dma_mm_read_read
	wire    [3:0] video_dma_mm_read_byteenable;                                                 // video_dma:mm_read_byteenable -> mm_interconnect_1:video_dma_mm_read_byteenable
	wire          video_dma_mm_read_readdatavalid;                                              // mm_interconnect_1:video_dma_mm_read_readdatavalid -> video_dma:mm_read_readdatavalid
	wire    [7:0] video_dma_mm_read_burstcount;                                                 // video_dma:mm_read_burstcount -> mm_interconnect_1:video_dma_mm_read_burstcount
	wire   [31:0] mdma_to_idct_accel_mm_read_readdata;                                          // mm_interconnect_1:mdma_to_idct_accel_mm_read_readdata -> mdma_to_idct_accel:mm_read_readdata
	wire          mdma_to_idct_accel_mm_read_waitrequest;                                       // mm_interconnect_1:mdma_to_idct_accel_mm_read_waitrequest -> mdma_to_idct_accel:mm_read_waitrequest
	wire   [28:0] mdma_to_idct_accel_mm_read_address;                                           // mdma_to_idct_accel:mm_read_address -> mm_interconnect_1:mdma_to_idct_accel_mm_read_address
	wire          mdma_to_idct_accel_mm_read_read;                                              // mdma_to_idct_accel:mm_read_read -> mm_interconnect_1:mdma_to_idct_accel_mm_read_read
	wire    [3:0] mdma_to_idct_accel_mm_read_byteenable;                                        // mdma_to_idct_accel:mm_read_byteenable -> mm_interconnect_1:mdma_to_idct_accel_mm_read_byteenable
	wire          mdma_to_idct_accel_mm_read_readdatavalid;                                     // mm_interconnect_1:mdma_to_idct_accel_mm_read_readdatavalid -> mdma_to_idct_accel:mm_read_readdatavalid
	wire    [7:0] mdma_to_idct_accel_mm_read_burstcount;                                        // mdma_to_idct_accel:mm_read_burstcount -> mm_interconnect_1:mdma_to_idct_accel_mm_read_burstcount
	wire   [31:0] mdma_to_ycbcr_to_rgb_accel_cb_mm_read_readdata;                               // mm_interconnect_1:mdma_to_ycbcr_to_rgb_accel_cb_mm_read_readdata -> mdma_to_ycbcr_to_rgb_accel_cb:mm_read_readdata
	wire          mdma_to_ycbcr_to_rgb_accel_cb_mm_read_waitrequest;                            // mm_interconnect_1:mdma_to_ycbcr_to_rgb_accel_cb_mm_read_waitrequest -> mdma_to_ycbcr_to_rgb_accel_cb:mm_read_waitrequest
	wire   [28:0] mdma_to_ycbcr_to_rgb_accel_cb_mm_read_address;                                // mdma_to_ycbcr_to_rgb_accel_cb:mm_read_address -> mm_interconnect_1:mdma_to_ycbcr_to_rgb_accel_cb_mm_read_address
	wire          mdma_to_ycbcr_to_rgb_accel_cb_mm_read_read;                                   // mdma_to_ycbcr_to_rgb_accel_cb:mm_read_read -> mm_interconnect_1:mdma_to_ycbcr_to_rgb_accel_cb_mm_read_read
	wire    [3:0] mdma_to_ycbcr_to_rgb_accel_cb_mm_read_byteenable;                             // mdma_to_ycbcr_to_rgb_accel_cb:mm_read_byteenable -> mm_interconnect_1:mdma_to_ycbcr_to_rgb_accel_cb_mm_read_byteenable
	wire          mdma_to_ycbcr_to_rgb_accel_cb_mm_read_readdatavalid;                          // mm_interconnect_1:mdma_to_ycbcr_to_rgb_accel_cb_mm_read_readdatavalid -> mdma_to_ycbcr_to_rgb_accel_cb:mm_read_readdatavalid
	wire    [7:0] mdma_to_ycbcr_to_rgb_accel_cb_mm_read_burstcount;                             // mdma_to_ycbcr_to_rgb_accel_cb:mm_read_burstcount -> mm_interconnect_1:mdma_to_ycbcr_to_rgb_accel_cb_mm_read_burstcount
	wire   [31:0] mdma_to_ycbcr_to_rgb_accel_cr_mm_read_readdata;                               // mm_interconnect_1:mdma_to_ycbcr_to_rgb_accel_cr_mm_read_readdata -> mdma_to_ycbcr_to_rgb_accel_cr:mm_read_readdata
	wire          mdma_to_ycbcr_to_rgb_accel_cr_mm_read_waitrequest;                            // mm_interconnect_1:mdma_to_ycbcr_to_rgb_accel_cr_mm_read_waitrequest -> mdma_to_ycbcr_to_rgb_accel_cr:mm_read_waitrequest
	wire   [28:0] mdma_to_ycbcr_to_rgb_accel_cr_mm_read_address;                                // mdma_to_ycbcr_to_rgb_accel_cr:mm_read_address -> mm_interconnect_1:mdma_to_ycbcr_to_rgb_accel_cr_mm_read_address
	wire          mdma_to_ycbcr_to_rgb_accel_cr_mm_read_read;                                   // mdma_to_ycbcr_to_rgb_accel_cr:mm_read_read -> mm_interconnect_1:mdma_to_ycbcr_to_rgb_accel_cr_mm_read_read
	wire    [3:0] mdma_to_ycbcr_to_rgb_accel_cr_mm_read_byteenable;                             // mdma_to_ycbcr_to_rgb_accel_cr:mm_read_byteenable -> mm_interconnect_1:mdma_to_ycbcr_to_rgb_accel_cr_mm_read_byteenable
	wire          mdma_to_ycbcr_to_rgb_accel_cr_mm_read_readdatavalid;                          // mm_interconnect_1:mdma_to_ycbcr_to_rgb_accel_cr_mm_read_readdatavalid -> mdma_to_ycbcr_to_rgb_accel_cr:mm_read_readdatavalid
	wire    [7:0] mdma_to_ycbcr_to_rgb_accel_cr_mm_read_burstcount;                             // mdma_to_ycbcr_to_rgb_accel_cr:mm_read_burstcount -> mm_interconnect_1:mdma_to_ycbcr_to_rgb_accel_cr_mm_read_burstcount
	wire   [31:0] mdma_to_ycbcr_to_rgb_accel_y_mm_read_readdata;                                // mm_interconnect_1:mdma_to_ycbcr_to_rgb_accel_y_mm_read_readdata -> mdma_to_ycbcr_to_rgb_accel_y:mm_read_readdata
	wire          mdma_to_ycbcr_to_rgb_accel_y_mm_read_waitrequest;                             // mm_interconnect_1:mdma_to_ycbcr_to_rgb_accel_y_mm_read_waitrequest -> mdma_to_ycbcr_to_rgb_accel_y:mm_read_waitrequest
	wire   [28:0] mdma_to_ycbcr_to_rgb_accel_y_mm_read_address;                                 // mdma_to_ycbcr_to_rgb_accel_y:mm_read_address -> mm_interconnect_1:mdma_to_ycbcr_to_rgb_accel_y_mm_read_address
	wire          mdma_to_ycbcr_to_rgb_accel_y_mm_read_read;                                    // mdma_to_ycbcr_to_rgb_accel_y:mm_read_read -> mm_interconnect_1:mdma_to_ycbcr_to_rgb_accel_y_mm_read_read
	wire    [3:0] mdma_to_ycbcr_to_rgb_accel_y_mm_read_byteenable;                              // mdma_to_ycbcr_to_rgb_accel_y:mm_read_byteenable -> mm_interconnect_1:mdma_to_ycbcr_to_rgb_accel_y_mm_read_byteenable
	wire          mdma_to_ycbcr_to_rgb_accel_y_mm_read_readdatavalid;                           // mm_interconnect_1:mdma_to_ycbcr_to_rgb_accel_y_mm_read_readdatavalid -> mdma_to_ycbcr_to_rgb_accel_y:mm_read_readdatavalid
	wire    [7:0] mdma_to_ycbcr_to_rgb_accel_y_mm_read_burstcount;                              // mdma_to_ycbcr_to_rgb_accel_y:mm_read_burstcount -> mm_interconnect_1:mdma_to_ycbcr_to_rgb_accel_y_mm_read_burstcount
	wire          mm_interconnect_1_lpddr2_avl_1_beginbursttransfer;                            // mm_interconnect_1:lpddr2_avl_1_beginbursttransfer -> lpddr2:avl_burstbegin_1
	wire   [31:0] mm_interconnect_1_lpddr2_avl_1_readdata;                                      // lpddr2:avl_rdata_1 -> mm_interconnect_1:lpddr2_avl_1_readdata
	wire          mm_interconnect_1_lpddr2_avl_1_waitrequest;                                   // lpddr2:avl_ready_1 -> mm_interconnect_1:lpddr2_avl_1_waitrequest
	wire   [26:0] mm_interconnect_1_lpddr2_avl_1_address;                                       // mm_interconnect_1:lpddr2_avl_1_address -> lpddr2:avl_addr_1
	wire          mm_interconnect_1_lpddr2_avl_1_read;                                          // mm_interconnect_1:lpddr2_avl_1_read -> lpddr2:avl_read_req_1
	wire    [3:0] mm_interconnect_1_lpddr2_avl_1_byteenable;                                    // mm_interconnect_1:lpddr2_avl_1_byteenable -> lpddr2:avl_be_1
	wire          mm_interconnect_1_lpddr2_avl_1_readdatavalid;                                 // lpddr2:avl_rdata_valid_1 -> mm_interconnect_1:lpddr2_avl_1_readdatavalid
	wire          mm_interconnect_1_lpddr2_avl_1_write;                                         // mm_interconnect_1:lpddr2_avl_1_write -> lpddr2:avl_write_req_1
	wire   [31:0] mm_interconnect_1_lpddr2_avl_1_writedata;                                     // mm_interconnect_1:lpddr2_avl_1_writedata -> lpddr2:avl_wdata_1
	wire    [7:0] mm_interconnect_1_lpddr2_avl_1_burstcount;                                    // mm_interconnect_1:lpddr2_avl_1_burstcount -> lpddr2:avl_size_1
	wire          mdma_from_idct_accel_mm_write_waitrequest;                                    // mm_interconnect_2:mdma_from_idct_accel_mm_write_waitrequest -> mdma_from_idct_accel:mm_write_waitrequest
	wire   [28:0] mdma_from_idct_accel_mm_write_address;                                        // mdma_from_idct_accel:mm_write_address -> mm_interconnect_2:mdma_from_idct_accel_mm_write_address
	wire    [3:0] mdma_from_idct_accel_mm_write_byteenable;                                     // mdma_from_idct_accel:mm_write_byteenable -> mm_interconnect_2:mdma_from_idct_accel_mm_write_byteenable
	wire          mdma_from_idct_accel_mm_write_write;                                          // mdma_from_idct_accel:mm_write_write -> mm_interconnect_2:mdma_from_idct_accel_mm_write_write
	wire   [31:0] mdma_from_idct_accel_mm_write_writedata;                                      // mdma_from_idct_accel:mm_write_writedata -> mm_interconnect_2:mdma_from_idct_accel_mm_write_writedata
	wire    [7:0] mdma_from_idct_accel_mm_write_burstcount;                                     // mdma_from_idct_accel:mm_write_burstcount -> mm_interconnect_2:mdma_from_idct_accel_mm_write_burstcount
	wire          mdma_from_ycbcr_to_rgb_accel_mm_write_waitrequest;                            // mm_interconnect_2:mdma_from_ycbcr_to_rgb_accel_mm_write_waitrequest -> mdma_from_ycbcr_to_rgb_accel:mm_write_waitrequest
	wire   [28:0] mdma_from_ycbcr_to_rgb_accel_mm_write_address;                                // mdma_from_ycbcr_to_rgb_accel:mm_write_address -> mm_interconnect_2:mdma_from_ycbcr_to_rgb_accel_mm_write_address
	wire    [3:0] mdma_from_ycbcr_to_rgb_accel_mm_write_byteenable;                             // mdma_from_ycbcr_to_rgb_accel:mm_write_byteenable -> mm_interconnect_2:mdma_from_ycbcr_to_rgb_accel_mm_write_byteenable
	wire          mdma_from_ycbcr_to_rgb_accel_mm_write_write;                                  // mdma_from_ycbcr_to_rgb_accel:mm_write_write -> mm_interconnect_2:mdma_from_ycbcr_to_rgb_accel_mm_write_write
	wire   [31:0] mdma_from_ycbcr_to_rgb_accel_mm_write_writedata;                              // mdma_from_ycbcr_to_rgb_accel:mm_write_writedata -> mm_interconnect_2:mdma_from_ycbcr_to_rgb_accel_mm_write_writedata
	wire    [7:0] mdma_from_ycbcr_to_rgb_accel_mm_write_burstcount;                             // mdma_from_ycbcr_to_rgb_accel:mm_write_burstcount -> mm_interconnect_2:mdma_from_ycbcr_to_rgb_accel_mm_write_burstcount
	wire          mm_interconnect_2_lpddr2_avl_2_beginbursttransfer;                            // mm_interconnect_2:lpddr2_avl_2_beginbursttransfer -> lpddr2:avl_burstbegin_2
	wire   [31:0] mm_interconnect_2_lpddr2_avl_2_readdata;                                      // lpddr2:avl_rdata_2 -> mm_interconnect_2:lpddr2_avl_2_readdata
	wire          mm_interconnect_2_lpddr2_avl_2_waitrequest;                                   // lpddr2:avl_ready_2 -> mm_interconnect_2:lpddr2_avl_2_waitrequest
	wire   [26:0] mm_interconnect_2_lpddr2_avl_2_address;                                       // mm_interconnect_2:lpddr2_avl_2_address -> lpddr2:avl_addr_2
	wire          mm_interconnect_2_lpddr2_avl_2_read;                                          // mm_interconnect_2:lpddr2_avl_2_read -> lpddr2:avl_read_req_2
	wire    [3:0] mm_interconnect_2_lpddr2_avl_2_byteenable;                                    // mm_interconnect_2:lpddr2_avl_2_byteenable -> lpddr2:avl_be_2
	wire          mm_interconnect_2_lpddr2_avl_2_readdatavalid;                                 // lpddr2:avl_rdata_valid_2 -> mm_interconnect_2:lpddr2_avl_2_readdatavalid
	wire          mm_interconnect_2_lpddr2_avl_2_write;                                         // mm_interconnect_2:lpddr2_avl_2_write -> lpddr2:avl_write_req_2
	wire   [31:0] mm_interconnect_2_lpddr2_avl_2_writedata;                                     // mm_interconnect_2:lpddr2_avl_2_writedata -> lpddr2:avl_wdata_2
	wire    [7:0] mm_interconnect_2_lpddr2_avl_2_burstcount;                                    // mm_interconnect_2:lpddr2_avl_2_burstcount -> lpddr2:avl_size_2
	wire          irq_mapper_receiver0_irq;                                                     // video_dma:csr_irq_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                                     // mailbox_simple_cpu0_to_cpu1:irq_space -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                                     // mailbox_simple_cpu1_to_cpu0:irq_msg -> irq_mapper:receiver2_irq
	wire          irq_mapper_receiver3_irq;                                                     // timer_0_0:irq -> irq_mapper:receiver3_irq
	wire          irq_mapper_receiver4_irq;                                                     // jtag_uart_0:av_irq -> irq_mapper:receiver4_irq
	wire          irq_mapper_receiver5_irq;                                                     // key:irq -> irq_mapper:receiver5_irq
	wire          irq_mapper_receiver6_irq;                                                     // timer_0_1:irq -> irq_mapper:receiver6_irq
	wire   [31:0] cpu_0_irq_irq;                                                                // irq_mapper:sender_irq -> cpu_0:irq
	wire          irq_mapper_001_receiver0_irq;                                                 // mdma_to_idct_accel:csr_irq_irq -> irq_mapper_001:receiver0_irq
	wire          irq_mapper_001_receiver1_irq;                                                 // mdma_from_idct_accel:csr_irq_irq -> irq_mapper_001:receiver1_irq
	wire          irq_mapper_001_receiver2_irq;                                                 // mdma_from_ycbcr_to_rgb_accel:csr_irq_irq -> irq_mapper_001:receiver2_irq
	wire          irq_mapper_001_receiver3_irq;                                                 // mdma_to_ycbcr_to_rgb_accel_cb:csr_irq_irq -> irq_mapper_001:receiver3_irq
	wire          irq_mapper_001_receiver4_irq;                                                 // mdma_to_ycbcr_to_rgb_accel_cr:csr_irq_irq -> irq_mapper_001:receiver4_irq
	wire          irq_mapper_001_receiver5_irq;                                                 // mdma_to_ycbcr_to_rgb_accel_y:csr_irq_irq -> irq_mapper_001:receiver5_irq
	wire          irq_mapper_001_receiver6_irq;                                                 // mailbox_simple_cpu1_to_cpu0:irq_space -> irq_mapper_001:receiver6_irq
	wire          irq_mapper_001_receiver7_irq;                                                 // mailbox_simple_cpu0_to_cpu1:irq_msg -> irq_mapper_001:receiver7_irq
	wire          irq_mapper_001_receiver8_irq;                                                 // jtag_uart_1:av_irq -> irq_mapper_001:receiver8_irq
	wire          irq_mapper_001_receiver9_irq;                                                 // timer_1_1:irq -> irq_mapper_001:receiver9_irq
	wire          irq_mapper_001_receiver10_irq;                                                // timer_1_0:irq -> irq_mapper_001:receiver10_irq
	wire   [31:0] cpu_1_irq_irq;                                                                // irq_mapper_001:sender_irq -> cpu_1:irq
	wire          video_fifo_out_valid;                                                         // video_fifo:avalonst_source_valid -> avalon_st_adapter:in_0_valid
	wire   [31:0] video_fifo_out_data;                                                          // video_fifo:avalonst_source_data -> avalon_st_adapter:in_0_data
	wire          video_fifo_out_ready;                                                         // avalon_st_adapter:in_0_ready -> video_fifo:avalonst_source_ready
	wire          video_fifo_out_startofpacket;                                                 // video_fifo:avalonst_source_startofpacket -> avalon_st_adapter:in_0_startofpacket
	wire          video_fifo_out_endofpacket;                                                   // video_fifo:avalonst_source_endofpacket -> avalon_st_adapter:in_0_endofpacket
	wire    [1:0] video_fifo_out_empty;                                                         // video_fifo:avalonst_source_empty -> avalon_st_adapter:in_0_empty
	wire          avalon_st_adapter_out_0_valid;                                                // avalon_st_adapter:out_0_valid -> pixel_conv:valid_in
	wire   [31:0] avalon_st_adapter_out_0_data;                                                 // avalon_st_adapter:out_0_data -> pixel_conv:data_in
	wire          avalon_st_adapter_out_0_ready;                                                // pixel_conv:ready_out -> avalon_st_adapter:out_0_ready
	wire          avalon_st_adapter_out_0_startofpacket;                                        // avalon_st_adapter:out_0_startofpacket -> pixel_conv:sop_in
	wire          avalon_st_adapter_out_0_endofpacket;                                          // avalon_st_adapter:out_0_endofpacket -> pixel_conv:eop_in
	wire    [1:0] avalon_st_adapter_out_0_empty;                                                // avalon_st_adapter:out_0_empty -> pixel_conv:empty_in
	wire          video_dma_st_source_valid;                                                    // video_dma:st_source_valid -> avalon_st_adapter_001:in_0_valid
	wire   [31:0] video_dma_st_source_data;                                                     // video_dma:st_source_data -> avalon_st_adapter_001:in_0_data
	wire          video_dma_st_source_ready;                                                    // avalon_st_adapter_001:in_0_ready -> video_dma:st_source_ready
	wire          video_dma_st_source_startofpacket;                                            // video_dma:st_source_startofpacket -> avalon_st_adapter_001:in_0_startofpacket
	wire          video_dma_st_source_endofpacket;                                              // video_dma:st_source_endofpacket -> avalon_st_adapter_001:in_0_endofpacket
	wire    [1:0] video_dma_st_source_empty;                                                    // video_dma:st_source_empty -> avalon_st_adapter_001:in_0_empty
	wire          avalon_st_adapter_001_out_0_valid;                                            // avalon_st_adapter_001:out_0_valid -> video_fifo:avalonst_sink_valid
	wire   [31:0] avalon_st_adapter_001_out_0_data;                                             // avalon_st_adapter_001:out_0_data -> video_fifo:avalonst_sink_data
	wire          avalon_st_adapter_001_out_0_ready;                                            // video_fifo:avalonst_sink_ready -> avalon_st_adapter_001:out_0_ready
	wire          avalon_st_adapter_001_out_0_startofpacket;                                    // avalon_st_adapter_001:out_0_startofpacket -> video_fifo:avalonst_sink_startofpacket
	wire          avalon_st_adapter_001_out_0_endofpacket;                                      // avalon_st_adapter_001:out_0_endofpacket -> video_fifo:avalonst_sink_endofpacket
	wire    [1:0] avalon_st_adapter_001_out_0_empty;                                            // avalon_st_adapter_001:out_0_empty -> video_fifo:avalonst_sink_empty
	wire          rst_controller_reset_out_reset;                                               // rst_controller:reset_out -> [cpu_0:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:cpu_0_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire          rst_controller_reset_out_reset_req;                                           // rst_controller:reset_req -> [cpu_0:reset_req, rst_translator:reset_req_in]
	wire          cpu_0_debug_reset_request_reset;                                              // cpu_0:debug_reset_request -> rst_controller:reset_in0
	wire          rst_controller_001_reset_out_reset;                                           // rst_controller_001:reset_out -> [cpu_1:reset_n, irq_mapper_001:reset, jtag_uart_1:rst_n, mm_interconnect_0:cpu_1_reset_reset_bridge_in_reset_reset, rst_translator_001:in_reset]
	wire          rst_controller_001_reset_out_reset_req;                                       // rst_controller_001:reset_req -> [cpu_1:reset_req, rst_translator_001:reset_req_in]
	wire          cpu_1_debug_reset_request_reset;                                              // cpu_1:debug_reset_request -> rst_controller_001:reset_in0
	wire          rst_controller_002_reset_out_reset;                                           // rst_controller_002:reset_out -> [avalon_st_adapter:in_rst_0_reset, pixel_conv:reset_n, video:reset_n, video_fifo:rdreset_n]
	wire          rst_controller_003_reset_out_reset;                                           // rst_controller_003:reset_out -> [mm_interconnect_0:sd_cont_reset_reset_bridge_in_reset_reset, sd_cont:reset]

	ECE423_QSYS_cpu_0 cpu_0 (
		.clk                                 (clk_125_clk),                                         //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (cpu_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_0_data_master_read),                              //                          .read
		.d_readdata                          (cpu_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_0_data_master_write),                             //                          .write
		.d_writedata                         (cpu_0_data_master_writedata),                         //                          .writedata
		.d_burstcount                        (cpu_0_data_master_burstcount),                        //                          .burstcount
		.d_readdatavalid                     (cpu_0_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_0_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                     // custom_instruction_master.readra
	);

	ECE423_QSYS_cpu_1 cpu_1 (
		.clk                                 (clk_125_clk),                                         //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                 //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),              //                          .reset_req
		.d_address                           (cpu_1_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_1_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_1_data_master_read),                              //                          .read
		.d_readdata                          (cpu_1_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_1_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_1_data_master_write),                             //                          .write
		.d_writedata                         (cpu_1_data_master_writedata),                         //                          .writedata
		.d_burstcount                        (cpu_1_data_master_burstcount),                        //                          .burstcount
		.d_readdatavalid                     (cpu_1_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_1_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_1_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_1_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_1_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_1_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_1_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_1_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_1_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_1_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_1_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_1_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_1_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_1_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_1_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_1_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_1_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                     // custom_instruction_master.readra
	);

	ECE423_QSYS_i2c_scl i2c_scl (
		.clk        (clk_125_clk),                             //                 clk.clk
		.reset_n    (~reset_controller_0_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_i2c_scl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_i2c_scl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_i2c_scl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_i2c_scl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_i2c_scl_s1_readdata),   //                    .readdata
		.out_port   (i2c_scl_export)                           // external_connection.export
	);

	ECE423_QSYS_i2c_sda i2c_sda (
		.clk        (clk_125_clk),                             //                 clk.clk
		.reset_n    (~reset_controller_0_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_i2c_sda_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_i2c_sda_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_i2c_sda_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_i2c_sda_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_i2c_sda_s1_readdata),   //                    .readdata
		.bidir_port (i2c_sda_export)                           // external_connection.export
	);

	idct_2D_streaming_interface idct_accelerator_2d (
		.clk     (clk_125_clk),                                       //                   clock.clk
		.i_data  (mdma_to_idct_accel_st_source_data),                 //   avalon_streaming_sink.data
		.i_valid (mdma_to_idct_accel_st_source_valid),                //                        .valid
		.o_ready (mdma_to_idct_accel_st_source_ready),                //                        .ready
		.i_ready (idct_accelerator_2d_avalon_streaming_source_ready), // avalon_streaming_source.ready
		.o_data  (idct_accelerator_2d_avalon_streaming_source_data),  //                        .data
		.o_valid (idct_accelerator_2d_avalon_streaming_source_valid), //                        .valid
		.reset_n (~reset_controller_0_reset_out_reset)                //                 reset_n.reset_n
	);

	ECE423_QSYS_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_125_clk),                                                 //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver4_irq)                                     //               irq.irq
	);

	ECE423_QSYS_jtag_uart_0 jtag_uart_1 (
		.clk            (clk_125_clk),                                                 //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_001_receiver8_irq)                                 //               irq.irq
	);

	ECE423_QSYS_key key (
		.clk        (clk_125_clk),                         //                 clk.clk
		.reset_n    (~reset_controller_0_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_0_key_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_key_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_key_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_key_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_key_s1_readdata),   //                    .readdata
		.in_port    (key_export),                          // external_connection.export
		.irq        (irq_mapper_receiver5_irq)             //                 irq.irq
	);

	ECE423_QSYS_ledg ledg (
		.clk        (clk_125_clk),                          //                 clk.clk
		.reset_n    (~reset_controller_0_reset_out_reset),  //               reset.reset_n
		.address    (mm_interconnect_0_ledg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledg_s1_readdata),   //                    .readdata
		.out_port   (ledg_export)                           // external_connection.export
	);

	ECE423_QSYS_ledg ledr (
		.clk        (clk_125_clk),                          //                 clk.clk
		.reset_n    (~reset_controller_0_reset_out_reset),  //               reset.reset_n
		.address    (mm_interconnect_0_ledr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledr_s1_readdata),   //                    .readdata
		.out_port   (ledr_export)                           // external_connection.export
	);

	ECE423_QSYS_lpddr2 lpddr2 (
		.pll_ref_clk                (lpddr2_pll_ref_clk_clk),                            //        pll_ref_clk.clk
		.global_reset_n             (lpddr2_global_reset_reset_n),                       //       global_reset.reset_n
		.soft_reset_n               (~reset_controller_0_reset_out_reset),               //         soft_reset.reset_n
		.afi_clk                    (),                                                  //            afi_clk.clk
		.afi_half_clk               (),                                                  //       afi_half_clk.clk
		.afi_reset_n                (),                                                  //          afi_reset.reset_n
		.afi_reset_export_n         (),                                                  //   afi_reset_export.reset_n
		.mem_ca                     (lpddr2_mem_ca),                                     //             memory.mem_ca
		.mem_ck                     (lpddr2_mem_ck),                                     //                   .mem_ck
		.mem_ck_n                   (lpddr2_mem_ck_n),                                   //                   .mem_ck_n
		.mem_cke                    (lpddr2_mem_cke),                                    //                   .mem_cke
		.mem_cs_n                   (lpddr2_mem_cs_n),                                   //                   .mem_cs_n
		.mem_dm                     (lpddr2_mem_dm),                                     //                   .mem_dm
		.mem_dq                     (lpddr2_mem_dq),                                     //                   .mem_dq
		.mem_dqs                    (lpddr2_mem_dqs),                                    //                   .mem_dqs
		.mem_dqs_n                  (lpddr2_mem_dqs_n),                                  //                   .mem_dqs_n
		.avl_ready_0                (mm_interconnect_0_lpddr2_avl_0_waitrequest),        //              avl_0.waitrequest_n
		.avl_burstbegin_0           (mm_interconnect_0_lpddr2_avl_0_beginbursttransfer), //                   .beginbursttransfer
		.avl_addr_0                 (mm_interconnect_0_lpddr2_avl_0_address),            //                   .address
		.avl_rdata_valid_0          (mm_interconnect_0_lpddr2_avl_0_readdatavalid),      //                   .readdatavalid
		.avl_rdata_0                (mm_interconnect_0_lpddr2_avl_0_readdata),           //                   .readdata
		.avl_wdata_0                (mm_interconnect_0_lpddr2_avl_0_writedata),          //                   .writedata
		.avl_be_0                   (mm_interconnect_0_lpddr2_avl_0_byteenable),         //                   .byteenable
		.avl_read_req_0             (mm_interconnect_0_lpddr2_avl_0_read),               //                   .read
		.avl_write_req_0            (mm_interconnect_0_lpddr2_avl_0_write),              //                   .write
		.avl_size_0                 (mm_interconnect_0_lpddr2_avl_0_burstcount),         //                   .burstcount
		.avl_ready_1                (mm_interconnect_1_lpddr2_avl_1_waitrequest),        //              avl_1.waitrequest_n
		.avl_burstbegin_1           (mm_interconnect_1_lpddr2_avl_1_beginbursttransfer), //                   .beginbursttransfer
		.avl_addr_1                 (mm_interconnect_1_lpddr2_avl_1_address),            //                   .address
		.avl_rdata_valid_1          (mm_interconnect_1_lpddr2_avl_1_readdatavalid),      //                   .readdatavalid
		.avl_rdata_1                (mm_interconnect_1_lpddr2_avl_1_readdata),           //                   .readdata
		.avl_wdata_1                (mm_interconnect_1_lpddr2_avl_1_writedata),          //                   .writedata
		.avl_be_1                   (mm_interconnect_1_lpddr2_avl_1_byteenable),         //                   .byteenable
		.avl_read_req_1             (mm_interconnect_1_lpddr2_avl_1_read),               //                   .read
		.avl_write_req_1            (mm_interconnect_1_lpddr2_avl_1_write),              //                   .write
		.avl_size_1                 (mm_interconnect_1_lpddr2_avl_1_burstcount),         //                   .burstcount
		.avl_ready_2                (mm_interconnect_2_lpddr2_avl_2_waitrequest),        //              avl_2.waitrequest_n
		.avl_burstbegin_2           (mm_interconnect_2_lpddr2_avl_2_beginbursttransfer), //                   .beginbursttransfer
		.avl_addr_2                 (mm_interconnect_2_lpddr2_avl_2_address),            //                   .address
		.avl_rdata_valid_2          (mm_interconnect_2_lpddr2_avl_2_readdatavalid),      //                   .readdatavalid
		.avl_rdata_2                (mm_interconnect_2_lpddr2_avl_2_readdata),           //                   .readdata
		.avl_wdata_2                (mm_interconnect_2_lpddr2_avl_2_writedata),          //                   .writedata
		.avl_be_2                   (mm_interconnect_2_lpddr2_avl_2_byteenable),         //                   .byteenable
		.avl_read_req_2             (mm_interconnect_2_lpddr2_avl_2_read),               //                   .read
		.avl_write_req_2            (mm_interconnect_2_lpddr2_avl_2_write),              //                   .write
		.avl_size_2                 (mm_interconnect_2_lpddr2_avl_2_burstcount),         //                   .burstcount
		.mp_cmd_clk_0_clk           (clk_125_clk),                                       //       mp_cmd_clk_0.clk
		.mp_cmd_reset_n_0_reset_n   (~reset_controller_0_reset_out_reset),               //   mp_cmd_reset_n_0.reset_n
		.mp_cmd_clk_1_clk           (clk_125_clk),                                       //       mp_cmd_clk_1.clk
		.mp_cmd_reset_n_1_reset_n   (~reset_controller_0_reset_out_reset),               //   mp_cmd_reset_n_1.reset_n
		.mp_cmd_clk_2_clk           (clk_125_clk),                                       //       mp_cmd_clk_2.clk
		.mp_cmd_reset_n_2_reset_n   (~reset_controller_0_reset_out_reset),               //   mp_cmd_reset_n_2.reset_n
		.mp_rfifo_clk_0_clk         (clk_125_clk),                                       //     mp_rfifo_clk_0.clk
		.mp_rfifo_reset_n_0_reset_n (~reset_controller_0_reset_out_reset),               // mp_rfifo_reset_n_0.reset_n
		.mp_wfifo_clk_0_clk         (clk_125_clk),                                       //     mp_wfifo_clk_0.clk
		.mp_wfifo_reset_n_0_reset_n (~reset_controller_0_reset_out_reset),               // mp_wfifo_reset_n_0.reset_n
		.mp_rfifo_clk_1_clk         (clk_125_clk),                                       //     mp_rfifo_clk_1.clk
		.mp_rfifo_reset_n_1_reset_n (~reset_controller_0_reset_out_reset),               // mp_rfifo_reset_n_1.reset_n
		.mp_wfifo_clk_1_clk         (clk_125_clk),                                       //     mp_wfifo_clk_1.clk
		.mp_wfifo_reset_n_1_reset_n (~reset_controller_0_reset_out_reset),               // mp_wfifo_reset_n_1.reset_n
		.local_init_done            (lpddr2_status_local_init_done),                     //             status.local_init_done
		.local_cal_success          (lpddr2_status_local_cal_success),                   //                   .local_cal_success
		.local_cal_fail             (lpddr2_status_local_cal_fail),                      //                   .local_cal_fail
		.oct_rzqin                  (lpddr2_oct_rzqin),                                  //                oct.rzqin
		.pll_mem_clk                (lpddr2_pll_sharing_pll_mem_clk),                    //        pll_sharing.pll_mem_clk
		.pll_write_clk              (lpddr2_pll_sharing_pll_write_clk),                  //                   .pll_write_clk
		.pll_locked                 (lpddr2_pll_sharing_pll_locked),                     //                   .pll_locked
		.pll_write_clk_pre_phy_clk  (lpddr2_pll_sharing_pll_write_clk_pre_phy_clk),      //                   .pll_write_clk_pre_phy_clk
		.pll_addr_cmd_clk           (lpddr2_pll_sharing_pll_addr_cmd_clk),               //                   .pll_addr_cmd_clk
		.pll_avl_clk                (lpddr2_pll_sharing_pll_avl_clk),                    //                   .pll_avl_clk
		.pll_config_clk             (lpddr2_pll_sharing_pll_config_clk),                 //                   .pll_config_clk
		.pll_mem_phy_clk            (lpddr2_pll_sharing_pll_mem_phy_clk),                //                   .pll_mem_phy_clk
		.afi_phy_clk                (lpddr2_pll_sharing_afi_phy_clk),                    //                   .afi_phy_clk
		.pll_avl_phy_clk            (lpddr2_pll_sharing_pll_avl_phy_clk)                 //                   .pll_avl_phy_clk
	);

	altera_avalon_mailbox #(
		.DWIDTH (32),
		.AWIDTH (2)
	) mailbox_simple_cpu0_to_cpu1 (
		.clk                  (clk_125_clk),                                                               //                    clk.clk
		.rst_n                (~reset_controller_0_reset_out_reset),                                       //                  rst_n.reset_n
		.avmm_snd_address     (mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_sender_address),     //        avmm_msg_sender.address
		.avmm_snd_writedata   (mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_sender_writedata),   //                       .writedata
		.avmm_snd_write       (mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_sender_write),       //                       .write
		.avmm_snd_read        (mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_sender_read),        //                       .read
		.avmm_snd_readdata    (mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_sender_readdata),    //                       .readdata
		.avmm_snd_waitrequest (mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_sender_waitrequest), //                       .waitrequest
		.irq_space            (irq_mapper_receiver1_irq),                                                  // interrupt_mb_available.irq
		.irq_msg              (irq_mapper_001_receiver7_irq),                                              //  interrupt_msg_pending.irq
		.avmm_rcv_address     (mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_receiver_address),   //      avmm_msg_receiver.address
		.avmm_rcv_read        (mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_receiver_read),      //                       .read
		.avmm_rcv_writedata   (mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_receiver_writedata), //                       .writedata
		.avmm_rcv_write       (mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_receiver_write),     //                       .write
		.avmm_rcv_readdata    (mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_receiver_readdata)   //                       .readdata
	);

	altera_avalon_mailbox #(
		.DWIDTH (32),
		.AWIDTH (2)
	) mailbox_simple_cpu1_to_cpu0 (
		.clk                  (clk_125_clk),                                                               //                    clk.clk
		.rst_n                (~reset_controller_0_reset_out_reset),                                       //                  rst_n.reset_n
		.avmm_snd_address     (mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_sender_address),     //        avmm_msg_sender.address
		.avmm_snd_writedata   (mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_sender_writedata),   //                       .writedata
		.avmm_snd_write       (mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_sender_write),       //                       .write
		.avmm_snd_read        (mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_sender_read),        //                       .read
		.avmm_snd_readdata    (mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_sender_readdata),    //                       .readdata
		.avmm_snd_waitrequest (mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_sender_waitrequest), //                       .waitrequest
		.irq_space            (irq_mapper_001_receiver6_irq),                                              // interrupt_mb_available.irq
		.irq_msg              (irq_mapper_receiver2_irq),                                                  //  interrupt_msg_pending.irq
		.avmm_rcv_address     (mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_receiver_address),   //      avmm_msg_receiver.address
		.avmm_rcv_read        (mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_receiver_read),      //                       .read
		.avmm_rcv_writedata   (mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_receiver_writedata), //                       .writedata
		.avmm_rcv_write       (mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_receiver_write),     //                       .write
		.avmm_rcv_readdata    (mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_receiver_readdata)   //                       .readdata
	);

	ECE423_QSYS_mdma_from_idct_accel mdma_from_idct_accel (
		.mm_write_address             (mdma_from_idct_accel_mm_write_address),                               //         mm_write.address
		.mm_write_write               (mdma_from_idct_accel_mm_write_write),                                 //                 .write
		.mm_write_byteenable          (mdma_from_idct_accel_mm_write_byteenable),                            //                 .byteenable
		.mm_write_writedata           (mdma_from_idct_accel_mm_write_writedata),                             //                 .writedata
		.mm_write_waitrequest         (mdma_from_idct_accel_mm_write_waitrequest),                           //                 .waitrequest
		.mm_write_burstcount          (mdma_from_idct_accel_mm_write_burstcount),                            //                 .burstcount
		.clock_clk                    (clk_125_clk),                                                         //            clock.clk
		.reset_n_reset_n              (~reset_controller_0_reset_out_reset),                                 //          reset_n.reset_n
		.csr_writedata                (mm_interconnect_0_mdma_from_idct_accel_csr_writedata),                //              csr.writedata
		.csr_write                    (mm_interconnect_0_mdma_from_idct_accel_csr_write),                    //                 .write
		.csr_byteenable               (mm_interconnect_0_mdma_from_idct_accel_csr_byteenable),               //                 .byteenable
		.csr_readdata                 (mm_interconnect_0_mdma_from_idct_accel_csr_readdata),                 //                 .readdata
		.csr_read                     (mm_interconnect_0_mdma_from_idct_accel_csr_read),                     //                 .read
		.csr_address                  (mm_interconnect_0_mdma_from_idct_accel_csr_address),                  //                 .address
		.descriptor_slave_write       (mm_interconnect_0_mdma_from_idct_accel_descriptor_slave_write),       // descriptor_slave.write
		.descriptor_slave_waitrequest (mm_interconnect_0_mdma_from_idct_accel_descriptor_slave_waitrequest), //                 .waitrequest
		.descriptor_slave_writedata   (mm_interconnect_0_mdma_from_idct_accel_descriptor_slave_writedata),   //                 .writedata
		.descriptor_slave_byteenable  (mm_interconnect_0_mdma_from_idct_accel_descriptor_slave_byteenable),  //                 .byteenable
		.csr_irq_irq                  (irq_mapper_001_receiver1_irq),                                        //          csr_irq.irq
		.st_sink_data                 (idct_accelerator_2d_avalon_streaming_source_data),                    //          st_sink.data
		.st_sink_valid                (idct_accelerator_2d_avalon_streaming_source_valid),                   //                 .valid
		.st_sink_ready                (idct_accelerator_2d_avalon_streaming_source_ready)                    //                 .ready
	);

	ECE423_QSYS_mdma_from_idct_accel mdma_from_ycbcr_to_rgb_accel (
		.mm_write_address             (mdma_from_ycbcr_to_rgb_accel_mm_write_address),                               //         mm_write.address
		.mm_write_write               (mdma_from_ycbcr_to_rgb_accel_mm_write_write),                                 //                 .write
		.mm_write_byteenable          (mdma_from_ycbcr_to_rgb_accel_mm_write_byteenable),                            //                 .byteenable
		.mm_write_writedata           (mdma_from_ycbcr_to_rgb_accel_mm_write_writedata),                             //                 .writedata
		.mm_write_waitrequest         (mdma_from_ycbcr_to_rgb_accel_mm_write_waitrequest),                           //                 .waitrequest
		.mm_write_burstcount          (mdma_from_ycbcr_to_rgb_accel_mm_write_burstcount),                            //                 .burstcount
		.clock_clk                    (clk_125_clk),                                                                 //            clock.clk
		.reset_n_reset_n              (~reset_controller_0_reset_out_reset),                                         //          reset_n.reset_n
		.csr_writedata                (mm_interconnect_0_mdma_from_ycbcr_to_rgb_accel_csr_writedata),                //              csr.writedata
		.csr_write                    (mm_interconnect_0_mdma_from_ycbcr_to_rgb_accel_csr_write),                    //                 .write
		.csr_byteenable               (mm_interconnect_0_mdma_from_ycbcr_to_rgb_accel_csr_byteenable),               //                 .byteenable
		.csr_readdata                 (mm_interconnect_0_mdma_from_ycbcr_to_rgb_accel_csr_readdata),                 //                 .readdata
		.csr_read                     (mm_interconnect_0_mdma_from_ycbcr_to_rgb_accel_csr_read),                     //                 .read
		.csr_address                  (mm_interconnect_0_mdma_from_ycbcr_to_rgb_accel_csr_address),                  //                 .address
		.descriptor_slave_write       (mm_interconnect_0_mdma_from_ycbcr_to_rgb_accel_descriptor_slave_write),       // descriptor_slave.write
		.descriptor_slave_waitrequest (mm_interconnect_0_mdma_from_ycbcr_to_rgb_accel_descriptor_slave_waitrequest), //                 .waitrequest
		.descriptor_slave_writedata   (mm_interconnect_0_mdma_from_ycbcr_to_rgb_accel_descriptor_slave_writedata),   //                 .writedata
		.descriptor_slave_byteenable  (mm_interconnect_0_mdma_from_ycbcr_to_rgb_accel_descriptor_slave_byteenable),  //                 .byteenable
		.csr_irq_irq                  (irq_mapper_001_receiver2_irq),                                                //          csr_irq.irq
		.st_sink_data                 (ycbcr_to_rgb_accelerator_avalon_streaming_source_data),                       //          st_sink.data
		.st_sink_valid                (ycbcr_to_rgb_accelerator_avalon_streaming_source_valid),                      //                 .valid
		.st_sink_ready                (ycbcr_to_rgb_accelerator_avalon_streaming_source_ready)                       //                 .ready
	);

	ECE423_QSYS_mdma_to_idct_accel mdma_to_idct_accel (
		.mm_read_address              (mdma_to_idct_accel_mm_read_address),                                //          mm_read.address
		.mm_read_read                 (mdma_to_idct_accel_mm_read_read),                                   //                 .read
		.mm_read_byteenable           (mdma_to_idct_accel_mm_read_byteenable),                             //                 .byteenable
		.mm_read_readdata             (mdma_to_idct_accel_mm_read_readdata),                               //                 .readdata
		.mm_read_waitrequest          (mdma_to_idct_accel_mm_read_waitrequest),                            //                 .waitrequest
		.mm_read_readdatavalid        (mdma_to_idct_accel_mm_read_readdatavalid),                          //                 .readdatavalid
		.mm_read_burstcount           (mdma_to_idct_accel_mm_read_burstcount),                             //                 .burstcount
		.clock_clk                    (clk_125_clk),                                                       //            clock.clk
		.reset_n_reset_n              (~reset_controller_0_reset_out_reset),                               //          reset_n.reset_n
		.csr_writedata                (mm_interconnect_0_mdma_to_idct_accel_csr_writedata),                //              csr.writedata
		.csr_write                    (mm_interconnect_0_mdma_to_idct_accel_csr_write),                    //                 .write
		.csr_byteenable               (mm_interconnect_0_mdma_to_idct_accel_csr_byteenable),               //                 .byteenable
		.csr_readdata                 (mm_interconnect_0_mdma_to_idct_accel_csr_readdata),                 //                 .readdata
		.csr_read                     (mm_interconnect_0_mdma_to_idct_accel_csr_read),                     //                 .read
		.csr_address                  (mm_interconnect_0_mdma_to_idct_accel_csr_address),                  //                 .address
		.descriptor_slave_write       (mm_interconnect_0_mdma_to_idct_accel_descriptor_slave_write),       // descriptor_slave.write
		.descriptor_slave_waitrequest (mm_interconnect_0_mdma_to_idct_accel_descriptor_slave_waitrequest), //                 .waitrequest
		.descriptor_slave_writedata   (mm_interconnect_0_mdma_to_idct_accel_descriptor_slave_writedata),   //                 .writedata
		.descriptor_slave_byteenable  (mm_interconnect_0_mdma_to_idct_accel_descriptor_slave_byteenable),  //                 .byteenable
		.csr_irq_irq                  (irq_mapper_001_receiver0_irq),                                      //          csr_irq.irq
		.st_source_data               (mdma_to_idct_accel_st_source_data),                                 //        st_source.data
		.st_source_valid              (mdma_to_idct_accel_st_source_valid),                                //                 .valid
		.st_source_ready              (mdma_to_idct_accel_st_source_ready)                                 //                 .ready
	);

	ECE423_QSYS_mdma_to_idct_accel mdma_to_ycbcr_to_rgb_accel_cb (
		.mm_read_address              (mdma_to_ycbcr_to_rgb_accel_cb_mm_read_address),                                //          mm_read.address
		.mm_read_read                 (mdma_to_ycbcr_to_rgb_accel_cb_mm_read_read),                                   //                 .read
		.mm_read_byteenable           (mdma_to_ycbcr_to_rgb_accel_cb_mm_read_byteenable),                             //                 .byteenable
		.mm_read_readdata             (mdma_to_ycbcr_to_rgb_accel_cb_mm_read_readdata),                               //                 .readdata
		.mm_read_waitrequest          (mdma_to_ycbcr_to_rgb_accel_cb_mm_read_waitrequest),                            //                 .waitrequest
		.mm_read_readdatavalid        (mdma_to_ycbcr_to_rgb_accel_cb_mm_read_readdatavalid),                          //                 .readdatavalid
		.mm_read_burstcount           (mdma_to_ycbcr_to_rgb_accel_cb_mm_read_burstcount),                             //                 .burstcount
		.clock_clk                    (clk_125_clk),                                                                  //            clock.clk
		.reset_n_reset_n              (~reset_controller_0_reset_out_reset),                                          //          reset_n.reset_n
		.csr_writedata                (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cb_csr_writedata),                //              csr.writedata
		.csr_write                    (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cb_csr_write),                    //                 .write
		.csr_byteenable               (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cb_csr_byteenable),               //                 .byteenable
		.csr_readdata                 (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cb_csr_readdata),                 //                 .readdata
		.csr_read                     (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cb_csr_read),                     //                 .read
		.csr_address                  (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cb_csr_address),                  //                 .address
		.descriptor_slave_write       (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cb_descriptor_slave_write),       // descriptor_slave.write
		.descriptor_slave_waitrequest (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cb_descriptor_slave_waitrequest), //                 .waitrequest
		.descriptor_slave_writedata   (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cb_descriptor_slave_writedata),   //                 .writedata
		.descriptor_slave_byteenable  (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cb_descriptor_slave_byteenable),  //                 .byteenable
		.csr_irq_irq                  (irq_mapper_001_receiver3_irq),                                                 //          csr_irq.irq
		.st_source_data               (mdma_to_ycbcr_to_rgb_accel_cb_st_source_data),                                 //        st_source.data
		.st_source_valid              (mdma_to_ycbcr_to_rgb_accel_cb_st_source_valid),                                //                 .valid
		.st_source_ready              (mdma_to_ycbcr_to_rgb_accel_cb_st_source_ready)                                 //                 .ready
	);

	ECE423_QSYS_mdma_to_idct_accel mdma_to_ycbcr_to_rgb_accel_cr (
		.mm_read_address              (mdma_to_ycbcr_to_rgb_accel_cr_mm_read_address),                                //          mm_read.address
		.mm_read_read                 (mdma_to_ycbcr_to_rgb_accel_cr_mm_read_read),                                   //                 .read
		.mm_read_byteenable           (mdma_to_ycbcr_to_rgb_accel_cr_mm_read_byteenable),                             //                 .byteenable
		.mm_read_readdata             (mdma_to_ycbcr_to_rgb_accel_cr_mm_read_readdata),                               //                 .readdata
		.mm_read_waitrequest          (mdma_to_ycbcr_to_rgb_accel_cr_mm_read_waitrequest),                            //                 .waitrequest
		.mm_read_readdatavalid        (mdma_to_ycbcr_to_rgb_accel_cr_mm_read_readdatavalid),                          //                 .readdatavalid
		.mm_read_burstcount           (mdma_to_ycbcr_to_rgb_accel_cr_mm_read_burstcount),                             //                 .burstcount
		.clock_clk                    (clk_125_clk),                                                                  //            clock.clk
		.reset_n_reset_n              (~reset_controller_0_reset_out_reset),                                          //          reset_n.reset_n
		.csr_writedata                (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cr_csr_writedata),                //              csr.writedata
		.csr_write                    (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cr_csr_write),                    //                 .write
		.csr_byteenable               (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cr_csr_byteenable),               //                 .byteenable
		.csr_readdata                 (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cr_csr_readdata),                 //                 .readdata
		.csr_read                     (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cr_csr_read),                     //                 .read
		.csr_address                  (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cr_csr_address),                  //                 .address
		.descriptor_slave_write       (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cr_descriptor_slave_write),       // descriptor_slave.write
		.descriptor_slave_waitrequest (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cr_descriptor_slave_waitrequest), //                 .waitrequest
		.descriptor_slave_writedata   (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cr_descriptor_slave_writedata),   //                 .writedata
		.descriptor_slave_byteenable  (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cr_descriptor_slave_byteenable),  //                 .byteenable
		.csr_irq_irq                  (irq_mapper_001_receiver4_irq),                                                 //          csr_irq.irq
		.st_source_data               (mdma_to_ycbcr_to_rgb_accel_cr_st_source_data),                                 //        st_source.data
		.st_source_valid              (mdma_to_ycbcr_to_rgb_accel_cr_st_source_valid),                                //                 .valid
		.st_source_ready              (mdma_to_ycbcr_to_rgb_accel_cr_st_source_ready)                                 //                 .ready
	);

	ECE423_QSYS_mdma_to_idct_accel mdma_to_ycbcr_to_rgb_accel_y (
		.mm_read_address              (mdma_to_ycbcr_to_rgb_accel_y_mm_read_address),                                //          mm_read.address
		.mm_read_read                 (mdma_to_ycbcr_to_rgb_accel_y_mm_read_read),                                   //                 .read
		.mm_read_byteenable           (mdma_to_ycbcr_to_rgb_accel_y_mm_read_byteenable),                             //                 .byteenable
		.mm_read_readdata             (mdma_to_ycbcr_to_rgb_accel_y_mm_read_readdata),                               //                 .readdata
		.mm_read_waitrequest          (mdma_to_ycbcr_to_rgb_accel_y_mm_read_waitrequest),                            //                 .waitrequest
		.mm_read_readdatavalid        (mdma_to_ycbcr_to_rgb_accel_y_mm_read_readdatavalid),                          //                 .readdatavalid
		.mm_read_burstcount           (mdma_to_ycbcr_to_rgb_accel_y_mm_read_burstcount),                             //                 .burstcount
		.clock_clk                    (clk_125_clk),                                                                 //            clock.clk
		.reset_n_reset_n              (~reset_controller_0_reset_out_reset),                                         //          reset_n.reset_n
		.csr_writedata                (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_y_csr_writedata),                //              csr.writedata
		.csr_write                    (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_y_csr_write),                    //                 .write
		.csr_byteenable               (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_y_csr_byteenable),               //                 .byteenable
		.csr_readdata                 (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_y_csr_readdata),                 //                 .readdata
		.csr_read                     (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_y_csr_read),                     //                 .read
		.csr_address                  (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_y_csr_address),                  //                 .address
		.descriptor_slave_write       (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_y_descriptor_slave_write),       // descriptor_slave.write
		.descriptor_slave_waitrequest (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_y_descriptor_slave_waitrequest), //                 .waitrequest
		.descriptor_slave_writedata   (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_y_descriptor_slave_writedata),   //                 .writedata
		.descriptor_slave_byteenable  (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_y_descriptor_slave_byteenable),  //                 .byteenable
		.csr_irq_irq                  (irq_mapper_001_receiver5_irq),                                                //          csr_irq.irq
		.st_source_data               (mdma_to_ycbcr_to_rgb_accel_y_st_source_data),                                 //        st_source.data
		.st_source_valid              (mdma_to_ycbcr_to_rgb_accel_y_st_source_valid),                                //                 .valid
		.st_source_ready              (mdma_to_ycbcr_to_rgb_accel_y_st_source_ready)                                 //                 .ready
	);

	ECE423_QSYS_mutex_0 mutex_0 (
		.reset_n       (~reset_controller_0_reset_out_reset),     // reset.reset_n
		.clk           (clk_125_clk),                             //   clk.clk
		.chipselect    (mm_interconnect_0_mutex_0_s1_chipselect), //    s1.chipselect
		.data_from_cpu (mm_interconnect_0_mutex_0_s1_writedata),  //      .writedata
		.read          (mm_interconnect_0_mutex_0_s1_read),       //      .read
		.write         (mm_interconnect_0_mutex_0_s1_write),      //      .write
		.data_to_cpu   (mm_interconnect_0_mutex_0_s1_readdata),   //      .readdata
		.address       (mm_interconnect_0_mutex_0_s1_address)     //      .address
	);

	Pixel_Conv #(
		.SOURCE_SYMBOLS_PER_BEAT (1)
	) pixel_conv (
		.clk       (video_clk_clk),                         //       clk.clk
		.reset_n   (~rst_controller_002_reset_out_reset),   // clk_reset.reset_n
		.ready_out (avalon_st_adapter_out_0_ready),         //        in.ready
		.valid_in  (avalon_st_adapter_out_0_valid),         //          .valid
		.data_in   (avalon_st_adapter_out_0_data),          //          .data
		.eop_in    (avalon_st_adapter_out_0_endofpacket),   //          .endofpacket
		.sop_in    (avalon_st_adapter_out_0_startofpacket), //          .startofpacket
		.empty_in  (avalon_st_adapter_out_0_empty),         //          .empty
		.ready_in  (pixel_conv_out_ready),                  //       out.ready
		.valid_out (pixel_conv_out_valid),                  //          .valid
		.data_out  (pixel_conv_out_data),                   //          .data
		.eop_out   (pixel_conv_out_endofpacket),            //          .endofpacket
		.sop_out   (pixel_conv_out_startofpacket),          //          .startofpacket
		.empty_out (pixel_conv_out_empty)                   //          .empty
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) reset_controller_0 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_125_clk),                        //       clk.clk
		.reset_out      (reset_controller_0_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	sd_cont sd_cont (
		.clk             (clk_50_clk),                                  //  clock.clk
		.reset           (rst_controller_003_reset_out_reset),          //  reset.reset
		.s_address       (mm_interconnect_0_sd_cont_slave_address),     //  slave.address
		.s_read          (mm_interconnect_0_sd_cont_slave_read),        //       .read
		.s_readdata      (mm_interconnect_0_sd_cont_slave_readdata),    //       .readdata
		.s_write         (mm_interconnect_0_sd_cont_slave_write),       //       .write
		.s_writedata     (mm_interconnect_0_sd_cont_slave_writedata),   //       .writedata
		.s_chipselect    (mm_interconnect_0_sd_cont_slave_chipselect),  //       .chipselect
		.s_waitrequest_n (mm_interconnect_0_sd_cont_slave_waitrequest), //       .waitrequest_n
		.m_address       (sd_cont_master_address),                      // master.address
		.m_read          (sd_cont_master_read),                         //       .read
		.m_readdata      (sd_cont_master_readdata),                     //       .readdata
		.m_write         (sd_cont_master_write),                        //       .write
		.m_writedata     (sd_cont_master_writedata),                    //       .writedata
		.m_waitrequest_n (~sd_cont_master_waitrequest),                 //       .waitrequest_n
		.sd_clk          (sd_sd_clk),                                   //     sd.sd_clk
		.sd_cmd          (sd_sd_cmd),                                   //       .sd_cmd
		.sd_dat          (sd_sd_dat),                                   //       .sd_dat
		.sd_pll_clk      (clk_50_clk)                                   // sd_clk.clk
	);

	ECE423_QSYS_sram #(
		.TCM_ADDRESS_W                  (19),
		.TCM_DATA_W                     (16),
		.TCM_BYTEENABLE_W               (2),
		.TCM_READ_WAIT                  (10),
		.TCM_WRITE_WAIT                 (10),
		.TCM_SETUP_WAIT                 (10),
		.TCM_DATA_HOLD                  (10),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (2),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (0),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (1),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (1),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (0),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (1),
		.ACTIVE_LOW_OUTPUTENABLE        (1),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) sram (
		.clk_clk                (clk_125_clk),                              //   clk.clk
		.reset_reset            (reset_controller_0_reset_out_reset),       // reset.reset
		.uas_address            (mm_interconnect_0_sram_uas_address),       //   uas.address
		.uas_burstcount         (mm_interconnect_0_sram_uas_burstcount),    //      .burstcount
		.uas_read               (mm_interconnect_0_sram_uas_read),          //      .read
		.uas_write              (mm_interconnect_0_sram_uas_write),         //      .write
		.uas_waitrequest        (mm_interconnect_0_sram_uas_waitrequest),   //      .waitrequest
		.uas_readdatavalid      (mm_interconnect_0_sram_uas_readdatavalid), //      .readdatavalid
		.uas_byteenable         (mm_interconnect_0_sram_uas_byteenable),    //      .byteenable
		.uas_readdata           (mm_interconnect_0_sram_uas_readdata),      //      .readdata
		.uas_writedata          (mm_interconnect_0_sram_uas_writedata),     //      .writedata
		.uas_lock               (mm_interconnect_0_sram_uas_lock),          //      .lock
		.uas_debugaccess        (mm_interconnect_0_sram_uas_debugaccess),   //      .debugaccess
		.tcm_write_n_out        (sram_tcm_write_n_out),                     //   tcm.write_n_out
		.tcm_chipselect_n_out   (sram_tcm_chipselect_n_out),                //      .chipselect_n_out
		.tcm_outputenable_n_out (sram_tcm_outputenable_n_out),              //      .outputenable_n_out
		.tcm_request            (sram_tcm_request),                         //      .request
		.tcm_grant              (sram_tcm_grant),                           //      .grant
		.tcm_address_out        (sram_tcm_address_out),                     //      .address_out
		.tcm_byteenable_n_out   (sram_tcm_byteenable_n_out),                //      .byteenable_n_out
		.tcm_data_out           (sram_tcm_data_out),                        //      .data_out
		.tcm_data_outen         (sram_tcm_data_outen),                      //      .data_outen
		.tcm_data_in            (sram_tcm_data_in)                          //      .data_in
	);

	ECE423_QSYS_sram_bridge sram_bridge (
		.clk                             (clk_125_clk),                                     //   clk.clk
		.reset                           (reset_controller_0_reset_out_reset),              // reset.reset
		.request                         (sram_sharer_tcm_request),                         //   tcs.request
		.grant                           (sram_sharer_tcm_grant),                           //      .grant
		.tcs_sram_tcm_data_out           (sram_sharer_tcm_sram_tcm_data_out_out),           //      .sram_tcm_data_out_out
		.tcs_sram_tcm_data_outen         (sram_sharer_tcm_sram_tcm_data_out_outen),         //      .sram_tcm_data_out_outen
		.tcs_sram_tcm_data_in            (sram_sharer_tcm_sram_tcm_data_out_in),            //      .sram_tcm_data_out_in
		.tcs_sram_tcm_address_out        (sram_sharer_tcm_sram_tcm_address_out_out),        //      .sram_tcm_address_out_out
		.tcs_sram_tcm_outputenable_n_out (sram_sharer_tcm_sram_tcm_outputenable_n_out_out), //      .sram_tcm_outputenable_n_out_out
		.tcs_sram_tcm_chipselect_n_out   (sram_sharer_tcm_sram_tcm_chipselect_n_out_out),   //      .sram_tcm_chipselect_n_out_out
		.tcs_sram_tcm_byteenable_n_out   (sram_sharer_tcm_sram_tcm_byteenable_n_out_out),   //      .sram_tcm_byteenable_n_out_out
		.tcs_sram_tcm_write_n_out        (sram_sharer_tcm_sram_tcm_write_n_out_out),        //      .sram_tcm_write_n_out_out
		.sram_tcm_data_out               (sram_bridge_out_sram_tcm_data_out),               //   out.sram_tcm_data_out
		.sram_tcm_address_out            (sram_bridge_out_sram_tcm_address_out),            //      .sram_tcm_address_out
		.sram_tcm_outputenable_n_out     (sram_bridge_out_sram_tcm_outputenable_n_out),     //      .sram_tcm_outputenable_n_out
		.sram_tcm_chipselect_n_out       (sram_bridge_out_sram_tcm_chipselect_n_out),       //      .sram_tcm_chipselect_n_out
		.sram_tcm_byteenable_n_out       (sram_bridge_out_sram_tcm_byteenable_n_out),       //      .sram_tcm_byteenable_n_out
		.sram_tcm_write_n_out            (sram_bridge_out_sram_tcm_write_n_out)             //      .sram_tcm_write_n_out
	);

	ECE423_QSYS_sram_sharer sram_sharer (
		.clk_clk                     (clk_125_clk),                                     //   clk.clk
		.reset_reset                 (reset_controller_0_reset_out_reset),              // reset.reset
		.request                     (sram_sharer_tcm_request),                         //   tcm.request
		.grant                       (sram_sharer_tcm_grant),                           //      .grant
		.sram_tcm_address_out        (sram_sharer_tcm_sram_tcm_address_out_out),        //      .sram_tcm_address_out_out
		.sram_tcm_byteenable_n_out   (sram_sharer_tcm_sram_tcm_byteenable_n_out_out),   //      .sram_tcm_byteenable_n_out_out
		.sram_tcm_outputenable_n_out (sram_sharer_tcm_sram_tcm_outputenable_n_out_out), //      .sram_tcm_outputenable_n_out_out
		.sram_tcm_write_n_out        (sram_sharer_tcm_sram_tcm_write_n_out_out),        //      .sram_tcm_write_n_out_out
		.sram_tcm_data_out           (sram_sharer_tcm_sram_tcm_data_out_out),           //      .sram_tcm_data_out_out
		.sram_tcm_data_in            (sram_sharer_tcm_sram_tcm_data_out_in),            //      .sram_tcm_data_out_in
		.sram_tcm_data_outen         (sram_sharer_tcm_sram_tcm_data_out_outen),         //      .sram_tcm_data_out_outen
		.sram_tcm_chipselect_n_out   (sram_sharer_tcm_sram_tcm_chipselect_n_out_out),   //      .sram_tcm_chipselect_n_out_out
		.tcs0_request                (sram_tcm_request),                                //  tcs0.request
		.tcs0_grant                  (sram_tcm_grant),                                  //      .grant
		.tcs0_address_out            (sram_tcm_address_out),                            //      .address_out
		.tcs0_byteenable_n_out       (sram_tcm_byteenable_n_out),                       //      .byteenable_n_out
		.tcs0_outputenable_n_out     (sram_tcm_outputenable_n_out),                     //      .outputenable_n_out
		.tcs0_write_n_out            (sram_tcm_write_n_out),                            //      .write_n_out
		.tcs0_data_out               (sram_tcm_data_out),                               //      .data_out
		.tcs0_data_in                (sram_tcm_data_in),                                //      .data_in
		.tcs0_data_outen             (sram_tcm_data_outen),                             //      .data_outen
		.tcs0_chipselect_n_out       (sram_tcm_chipselect_n_out)                        //      .chipselect_n_out
	);

	ECE423_QSYS_sysid sysid (
		.clock    (clk_125_clk),                                    //           clk.clk
		.reset_n  (~reset_controller_0_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	ECE423_QSYS_timer_0_0 timer_0_0 (
		.clk        (clk_125_clk),                               //   clk.clk
		.reset_n    (~reset_controller_0_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_0_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                   //   irq.irq
	);

	ECE423_QSYS_timer_0_1 timer_0_1 (
		.clk        (clk_125_clk),                               //   clk.clk
		.reset_n    (~reset_controller_0_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_0_1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_1_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver6_irq)                   //   irq.irq
	);

	ECE423_QSYS_timer_0_1 timer_1_0 (
		.clk        (clk_125_clk),                               //   clk.clk
		.reset_n    (~reset_controller_0_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_1_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1_0_s1_write),     //      .write_n
		.irq        (irq_mapper_001_receiver10_irq)              //   irq.irq
	);

	ECE423_QSYS_timer_0_1 timer_1_1 (
		.clk        (clk_125_clk),                               //   clk.clk
		.reset_n    (~reset_controller_0_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_1_1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1_1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1_1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1_1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1_1_s1_write),     //      .write_n
		.irq        (irq_mapper_001_receiver9_irq)               //   irq.irq
	);

	altera_avalon_video_sync_generator #(
		.DATA_STREAM_BIT_WIDTH (24),
		.BEATS_PER_PIXEL       (1),
		.NUM_COLUMNS           (640),
		.NUM_ROWS              (480),
		.H_BLANK_PIXELS        (128),
		.H_FRONT_PORCH_PIXELS  (24),
		.H_SYNC_PULSE_PIXELS   (32),
		.H_SYNC_PULSE_POLARITY (0),
		.V_BLANK_LINES         (45),
		.V_FRONT_PORCH_LINES   (10),
		.V_SYNC_PULSE_LINES    (3),
		.V_SYNC_PULSE_POLARITY (0),
		.TOTAL_HSCAN_PIXELS    (768),
		.TOTAL_VSCAN_LINES     (525)
	) video (
		.clk     (video_clk_clk),                       //       clk.clk
		.reset_n (~rst_controller_002_reset_out_reset), // clk_reset.reset_n
		.ready   (pixel_conv_out_ready),                //        in.ready
		.valid   (pixel_conv_out_valid),                //          .valid
		.data    (pixel_conv_out_data),                 //          .data
		.eop     (pixel_conv_out_endofpacket),          //          .endofpacket
		.sop     (pixel_conv_out_startofpacket),        //          .startofpacket
		.empty   (pixel_conv_out_empty),                //          .empty
		.RGB_OUT (video_RGB_OUT),                       //      sync.export
		.HD      (video_HD),                            //          .export
		.VD      (video_VD),                            //          .export
		.DEN     (video_DEN)                            //          .export
	);

	ECE423_QSYS_video_dma video_dma (
		.mm_read_address              (video_dma_mm_read_address),                                //          mm_read.address
		.mm_read_read                 (video_dma_mm_read_read),                                   //                 .read
		.mm_read_byteenable           (video_dma_mm_read_byteenable),                             //                 .byteenable
		.mm_read_readdata             (video_dma_mm_read_readdata),                               //                 .readdata
		.mm_read_waitrequest          (video_dma_mm_read_waitrequest),                            //                 .waitrequest
		.mm_read_readdatavalid        (video_dma_mm_read_readdatavalid),                          //                 .readdatavalid
		.mm_read_burstcount           (video_dma_mm_read_burstcount),                             //                 .burstcount
		.clock_clk                    (clk_125_clk),                                              //            clock.clk
		.reset_n_reset_n              (~reset_controller_0_reset_out_reset),                      //          reset_n.reset_n
		.csr_writedata                (mm_interconnect_0_video_dma_csr_writedata),                //              csr.writedata
		.csr_write                    (mm_interconnect_0_video_dma_csr_write),                    //                 .write
		.csr_byteenable               (mm_interconnect_0_video_dma_csr_byteenable),               //                 .byteenable
		.csr_readdata                 (mm_interconnect_0_video_dma_csr_readdata),                 //                 .readdata
		.csr_read                     (mm_interconnect_0_video_dma_csr_read),                     //                 .read
		.csr_address                  (mm_interconnect_0_video_dma_csr_address),                  //                 .address
		.descriptor_slave_write       (mm_interconnect_0_video_dma_descriptor_slave_write),       // descriptor_slave.write
		.descriptor_slave_waitrequest (mm_interconnect_0_video_dma_descriptor_slave_waitrequest), //                 .waitrequest
		.descriptor_slave_writedata   (mm_interconnect_0_video_dma_descriptor_slave_writedata),   //                 .writedata
		.descriptor_slave_byteenable  (mm_interconnect_0_video_dma_descriptor_slave_byteenable),  //                 .byteenable
		.csr_irq_irq                  (irq_mapper_receiver0_irq),                                 //          csr_irq.irq
		.st_source_data               (video_dma_st_source_data),                                 //        st_source.data
		.st_source_valid              (video_dma_st_source_valid),                                //                 .valid
		.st_source_ready              (video_dma_st_source_ready),                                //                 .ready
		.st_source_startofpacket      (video_dma_st_source_startofpacket),                        //                 .startofpacket
		.st_source_endofpacket        (video_dma_st_source_endofpacket),                          //                 .endofpacket
		.st_source_empty              (video_dma_st_source_empty)                                 //                 .empty
	);

	ECE423_QSYS_video_fifo video_fifo (
		.wrclock                       (clk_125_clk),                               //    clk_in.clk
		.wrreset_n                     (~reset_controller_0_reset_out_reset),       //  reset_in.reset_n
		.rdclock                       (video_clk_clk),                             //   clk_out.clk
		.rdreset_n                     (~rst_controller_002_reset_out_reset),       // reset_out.reset_n
		.avalonst_sink_valid           (avalon_st_adapter_001_out_0_valid),         //        in.valid
		.avalonst_sink_data            (avalon_st_adapter_001_out_0_data),          //          .data
		.avalonst_sink_startofpacket   (avalon_st_adapter_001_out_0_startofpacket), //          .startofpacket
		.avalonst_sink_endofpacket     (avalon_st_adapter_001_out_0_endofpacket),   //          .endofpacket
		.avalonst_sink_empty           (avalon_st_adapter_001_out_0_empty),         //          .empty
		.avalonst_sink_ready           (avalon_st_adapter_001_out_0_ready),         //          .ready
		.avalonst_source_valid         (video_fifo_out_valid),                      //       out.valid
		.avalonst_source_data          (video_fifo_out_data),                       //          .data
		.avalonst_source_startofpacket (video_fifo_out_startofpacket),              //          .startofpacket
		.avalonst_source_endofpacket   (video_fifo_out_endofpacket),                //          .endofpacket
		.avalonst_source_empty         (video_fifo_out_empty),                      //          .empty
		.avalonst_source_ready         (video_fifo_out_ready)                       //          .ready
	);

	ECE423_QSYS_video_pll video_pll (
		.refclk   (clk_50_clk),                         //  refclk.clk
		.rst      (reset_controller_0_reset_out_reset), //   reset.reset
		.outclk_0 (video_clk_clk),                      // outclk0.clk
		.locked   ()                                    // (terminated)
	);

	ycbcr_to_rgb_streaming_interface ycbcr_to_rgb_accelerator (
		.clk         (clk_125_clk),                                            //                    clock.clk
		.i_rgb_ready (ycbcr_to_rgb_accelerator_avalon_streaming_source_ready), //  avalon_streaming_source.ready
		.o_rgb_data  (ycbcr_to_rgb_accelerator_avalon_streaming_source_data),  //                         .data
		.o_rgb_valid (ycbcr_to_rgb_accelerator_avalon_streaming_source_valid), //                         .valid
		.o_cr_ready  (mdma_to_ycbcr_to_rgb_accel_cr_st_source_ready),          // avalon_streaming_sink_cr.ready
		.i_cr_data   (mdma_to_ycbcr_to_rgb_accel_cr_st_source_data),           //                         .data
		.i_cr_valid  (mdma_to_ycbcr_to_rgb_accel_cr_st_source_valid),          //                         .valid
		.o_y_ready   (mdma_to_ycbcr_to_rgb_accel_y_st_source_ready),           //  avalon_streaming_sink_y.ready
		.i_y_valid   (mdma_to_ycbcr_to_rgb_accel_y_st_source_valid),           //                         .valid
		.i_y_data    (mdma_to_ycbcr_to_rgb_accel_y_st_source_data),            //                         .data
		.i_cb_data   (mdma_to_ycbcr_to_rgb_accel_cb_st_source_data),           // avalon_streaming_sink_cb.data
		.i_cb_valid  (mdma_to_ycbcr_to_rgb_accel_cb_st_source_valid),          //                         .valid
		.o_cb_ready  (mdma_to_ycbcr_to_rgb_accel_cb_st_source_ready),          //                         .ready
		.reset_n     (~reset_controller_0_reset_out_reset)                     //                  reset_n.reset_n
	);

	ECE423_QSYS_mm_interconnect_0 mm_interconnect_0 (
		.clk_125_clk_clk                                               (clk_125_clk),                                                                  //                                             clk_125_clk.clk
		.clk_50_out_clk_clk                                            (clk_50_clk),                                                                   //                                          clk_50_out_clk.clk
		.cpu_0_reset_reset_bridge_in_reset_reset                       (rst_controller_reset_out_reset),                                               //                       cpu_0_reset_reset_bridge_in_reset.reset
		.cpu_1_reset_reset_bridge_in_reset_reset                       (rst_controller_001_reset_out_reset),                                           //                       cpu_1_reset_reset_bridge_in_reset.reset
		.lpddr2_mp_cmd_reset_n_0_reset_bridge_in_reset_reset           (reset_controller_0_reset_out_reset),                                           //           lpddr2_mp_cmd_reset_n_0_reset_bridge_in_reset.reset
		.mailbox_simple_cpu1_to_cpu0_rst_n_reset_bridge_in_reset_reset (reset_controller_0_reset_out_reset),                                           // mailbox_simple_cpu1_to_cpu0_rst_n_reset_bridge_in_reset.reset
		.sd_cont_reset_reset_bridge_in_reset_reset                     (rst_controller_003_reset_out_reset),                                           //                     sd_cont_reset_reset_bridge_in_reset.reset
		.cpu_0_data_master_address                                     (cpu_0_data_master_address),                                                    //                                       cpu_0_data_master.address
		.cpu_0_data_master_waitrequest                                 (cpu_0_data_master_waitrequest),                                                //                                                        .waitrequest
		.cpu_0_data_master_burstcount                                  (cpu_0_data_master_burstcount),                                                 //                                                        .burstcount
		.cpu_0_data_master_byteenable                                  (cpu_0_data_master_byteenable),                                                 //                                                        .byteenable
		.cpu_0_data_master_read                                        (cpu_0_data_master_read),                                                       //                                                        .read
		.cpu_0_data_master_readdata                                    (cpu_0_data_master_readdata),                                                   //                                                        .readdata
		.cpu_0_data_master_readdatavalid                               (cpu_0_data_master_readdatavalid),                                              //                                                        .readdatavalid
		.cpu_0_data_master_write                                       (cpu_0_data_master_write),                                                      //                                                        .write
		.cpu_0_data_master_writedata                                   (cpu_0_data_master_writedata),                                                  //                                                        .writedata
		.cpu_0_data_master_debugaccess                                 (cpu_0_data_master_debugaccess),                                                //                                                        .debugaccess
		.cpu_0_instruction_master_address                              (cpu_0_instruction_master_address),                                             //                                cpu_0_instruction_master.address
		.cpu_0_instruction_master_waitrequest                          (cpu_0_instruction_master_waitrequest),                                         //                                                        .waitrequest
		.cpu_0_instruction_master_read                                 (cpu_0_instruction_master_read),                                                //                                                        .read
		.cpu_0_instruction_master_readdata                             (cpu_0_instruction_master_readdata),                                            //                                                        .readdata
		.cpu_0_instruction_master_readdatavalid                        (cpu_0_instruction_master_readdatavalid),                                       //                                                        .readdatavalid
		.cpu_1_data_master_address                                     (cpu_1_data_master_address),                                                    //                                       cpu_1_data_master.address
		.cpu_1_data_master_waitrequest                                 (cpu_1_data_master_waitrequest),                                                //                                                        .waitrequest
		.cpu_1_data_master_burstcount                                  (cpu_1_data_master_burstcount),                                                 //                                                        .burstcount
		.cpu_1_data_master_byteenable                                  (cpu_1_data_master_byteenable),                                                 //                                                        .byteenable
		.cpu_1_data_master_read                                        (cpu_1_data_master_read),                                                       //                                                        .read
		.cpu_1_data_master_readdata                                    (cpu_1_data_master_readdata),                                                   //                                                        .readdata
		.cpu_1_data_master_readdatavalid                               (cpu_1_data_master_readdatavalid),                                              //                                                        .readdatavalid
		.cpu_1_data_master_write                                       (cpu_1_data_master_write),                                                      //                                                        .write
		.cpu_1_data_master_writedata                                   (cpu_1_data_master_writedata),                                                  //                                                        .writedata
		.cpu_1_data_master_debugaccess                                 (cpu_1_data_master_debugaccess),                                                //                                                        .debugaccess
		.cpu_1_instruction_master_address                              (cpu_1_instruction_master_address),                                             //                                cpu_1_instruction_master.address
		.cpu_1_instruction_master_waitrequest                          (cpu_1_instruction_master_waitrequest),                                         //                                                        .waitrequest
		.cpu_1_instruction_master_read                                 (cpu_1_instruction_master_read),                                                //                                                        .read
		.cpu_1_instruction_master_readdata                             (cpu_1_instruction_master_readdata),                                            //                                                        .readdata
		.cpu_1_instruction_master_readdatavalid                        (cpu_1_instruction_master_readdatavalid),                                       //                                                        .readdatavalid
		.sd_cont_master_address                                        (sd_cont_master_address),                                                       //                                          sd_cont_master.address
		.sd_cont_master_waitrequest                                    (sd_cont_master_waitrequest),                                                   //                                                        .waitrequest
		.sd_cont_master_read                                           (sd_cont_master_read),                                                          //                                                        .read
		.sd_cont_master_readdata                                       (sd_cont_master_readdata),                                                      //                                                        .readdata
		.sd_cont_master_write                                          (sd_cont_master_write),                                                         //                                                        .write
		.sd_cont_master_writedata                                      (sd_cont_master_writedata),                                                     //                                                        .writedata
		.cpu_0_debug_mem_slave_address                                 (mm_interconnect_0_cpu_0_debug_mem_slave_address),                              //                                   cpu_0_debug_mem_slave.address
		.cpu_0_debug_mem_slave_write                                   (mm_interconnect_0_cpu_0_debug_mem_slave_write),                                //                                                        .write
		.cpu_0_debug_mem_slave_read                                    (mm_interconnect_0_cpu_0_debug_mem_slave_read),                                 //                                                        .read
		.cpu_0_debug_mem_slave_readdata                                (mm_interconnect_0_cpu_0_debug_mem_slave_readdata),                             //                                                        .readdata
		.cpu_0_debug_mem_slave_writedata                               (mm_interconnect_0_cpu_0_debug_mem_slave_writedata),                            //                                                        .writedata
		.cpu_0_debug_mem_slave_byteenable                              (mm_interconnect_0_cpu_0_debug_mem_slave_byteenable),                           //                                                        .byteenable
		.cpu_0_debug_mem_slave_waitrequest                             (mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest),                          //                                                        .waitrequest
		.cpu_0_debug_mem_slave_debugaccess                             (mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess),                          //                                                        .debugaccess
		.cpu_1_debug_mem_slave_address                                 (mm_interconnect_0_cpu_1_debug_mem_slave_address),                              //                                   cpu_1_debug_mem_slave.address
		.cpu_1_debug_mem_slave_write                                   (mm_interconnect_0_cpu_1_debug_mem_slave_write),                                //                                                        .write
		.cpu_1_debug_mem_slave_read                                    (mm_interconnect_0_cpu_1_debug_mem_slave_read),                                 //                                                        .read
		.cpu_1_debug_mem_slave_readdata                                (mm_interconnect_0_cpu_1_debug_mem_slave_readdata),                             //                                                        .readdata
		.cpu_1_debug_mem_slave_writedata                               (mm_interconnect_0_cpu_1_debug_mem_slave_writedata),                            //                                                        .writedata
		.cpu_1_debug_mem_slave_byteenable                              (mm_interconnect_0_cpu_1_debug_mem_slave_byteenable),                           //                                                        .byteenable
		.cpu_1_debug_mem_slave_waitrequest                             (mm_interconnect_0_cpu_1_debug_mem_slave_waitrequest),                          //                                                        .waitrequest
		.cpu_1_debug_mem_slave_debugaccess                             (mm_interconnect_0_cpu_1_debug_mem_slave_debugaccess),                          //                                                        .debugaccess
		.i2c_scl_s1_address                                            (mm_interconnect_0_i2c_scl_s1_address),                                         //                                              i2c_scl_s1.address
		.i2c_scl_s1_write                                              (mm_interconnect_0_i2c_scl_s1_write),                                           //                                                        .write
		.i2c_scl_s1_readdata                                           (mm_interconnect_0_i2c_scl_s1_readdata),                                        //                                                        .readdata
		.i2c_scl_s1_writedata                                          (mm_interconnect_0_i2c_scl_s1_writedata),                                       //                                                        .writedata
		.i2c_scl_s1_chipselect                                         (mm_interconnect_0_i2c_scl_s1_chipselect),                                      //                                                        .chipselect
		.i2c_sda_s1_address                                            (mm_interconnect_0_i2c_sda_s1_address),                                         //                                              i2c_sda_s1.address
		.i2c_sda_s1_write                                              (mm_interconnect_0_i2c_sda_s1_write),                                           //                                                        .write
		.i2c_sda_s1_readdata                                           (mm_interconnect_0_i2c_sda_s1_readdata),                                        //                                                        .readdata
		.i2c_sda_s1_writedata                                          (mm_interconnect_0_i2c_sda_s1_writedata),                                       //                                                        .writedata
		.i2c_sda_s1_chipselect                                         (mm_interconnect_0_i2c_sda_s1_chipselect),                                      //                                                        .chipselect
		.jtag_uart_0_avalon_jtag_slave_address                         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),                      //                           jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),                        //                                                        .write
		.jtag_uart_0_avalon_jtag_slave_read                            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),                         //                                                        .read
		.jtag_uart_0_avalon_jtag_slave_readdata                        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),                     //                                                        .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),                    //                                                        .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),                  //                                                        .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),                   //                                                        .chipselect
		.jtag_uart_1_avalon_jtag_slave_address                         (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_address),                      //                           jtag_uart_1_avalon_jtag_slave.address
		.jtag_uart_1_avalon_jtag_slave_write                           (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write),                        //                                                        .write
		.jtag_uart_1_avalon_jtag_slave_read                            (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read),                         //                                                        .read
		.jtag_uart_1_avalon_jtag_slave_readdata                        (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_readdata),                     //                                                        .readdata
		.jtag_uart_1_avalon_jtag_slave_writedata                       (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_writedata),                    //                                                        .writedata
		.jtag_uart_1_avalon_jtag_slave_waitrequest                     (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_waitrequest),                  //                                                        .waitrequest
		.jtag_uart_1_avalon_jtag_slave_chipselect                      (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_chipselect),                   //                                                        .chipselect
		.key_s1_address                                                (mm_interconnect_0_key_s1_address),                                             //                                                  key_s1.address
		.key_s1_write                                                  (mm_interconnect_0_key_s1_write),                                               //                                                        .write
		.key_s1_readdata                                               (mm_interconnect_0_key_s1_readdata),                                            //                                                        .readdata
		.key_s1_writedata                                              (mm_interconnect_0_key_s1_writedata),                                           //                                                        .writedata
		.key_s1_chipselect                                             (mm_interconnect_0_key_s1_chipselect),                                          //                                                        .chipselect
		.ledg_s1_address                                               (mm_interconnect_0_ledg_s1_address),                                            //                                                 ledg_s1.address
		.ledg_s1_write                                                 (mm_interconnect_0_ledg_s1_write),                                              //                                                        .write
		.ledg_s1_readdata                                              (mm_interconnect_0_ledg_s1_readdata),                                           //                                                        .readdata
		.ledg_s1_writedata                                             (mm_interconnect_0_ledg_s1_writedata),                                          //                                                        .writedata
		.ledg_s1_chipselect                                            (mm_interconnect_0_ledg_s1_chipselect),                                         //                                                        .chipselect
		.ledr_s1_address                                               (mm_interconnect_0_ledr_s1_address),                                            //                                                 ledr_s1.address
		.ledr_s1_write                                                 (mm_interconnect_0_ledr_s1_write),                                              //                                                        .write
		.ledr_s1_readdata                                              (mm_interconnect_0_ledr_s1_readdata),                                           //                                                        .readdata
		.ledr_s1_writedata                                             (mm_interconnect_0_ledr_s1_writedata),                                          //                                                        .writedata
		.ledr_s1_chipselect                                            (mm_interconnect_0_ledr_s1_chipselect),                                         //                                                        .chipselect
		.lpddr2_avl_0_address                                          (mm_interconnect_0_lpddr2_avl_0_address),                                       //                                            lpddr2_avl_0.address
		.lpddr2_avl_0_write                                            (mm_interconnect_0_lpddr2_avl_0_write),                                         //                                                        .write
		.lpddr2_avl_0_read                                             (mm_interconnect_0_lpddr2_avl_0_read),                                          //                                                        .read
		.lpddr2_avl_0_readdata                                         (mm_interconnect_0_lpddr2_avl_0_readdata),                                      //                                                        .readdata
		.lpddr2_avl_0_writedata                                        (mm_interconnect_0_lpddr2_avl_0_writedata),                                     //                                                        .writedata
		.lpddr2_avl_0_beginbursttransfer                               (mm_interconnect_0_lpddr2_avl_0_beginbursttransfer),                            //                                                        .beginbursttransfer
		.lpddr2_avl_0_burstcount                                       (mm_interconnect_0_lpddr2_avl_0_burstcount),                                    //                                                        .burstcount
		.lpddr2_avl_0_byteenable                                       (mm_interconnect_0_lpddr2_avl_0_byteenable),                                    //                                                        .byteenable
		.lpddr2_avl_0_readdatavalid                                    (mm_interconnect_0_lpddr2_avl_0_readdatavalid),                                 //                                                        .readdatavalid
		.lpddr2_avl_0_waitrequest                                      (~mm_interconnect_0_lpddr2_avl_0_waitrequest),                                  //                                                        .waitrequest
		.mailbox_simple_cpu0_to_cpu1_avmm_msg_receiver_address         (mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_receiver_address),      //           mailbox_simple_cpu0_to_cpu1_avmm_msg_receiver.address
		.mailbox_simple_cpu0_to_cpu1_avmm_msg_receiver_write           (mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_receiver_write),        //                                                        .write
		.mailbox_simple_cpu0_to_cpu1_avmm_msg_receiver_read            (mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_receiver_read),         //                                                        .read
		.mailbox_simple_cpu0_to_cpu1_avmm_msg_receiver_readdata        (mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_receiver_readdata),     //                                                        .readdata
		.mailbox_simple_cpu0_to_cpu1_avmm_msg_receiver_writedata       (mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_receiver_writedata),    //                                                        .writedata
		.mailbox_simple_cpu0_to_cpu1_avmm_msg_sender_address           (mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_sender_address),        //             mailbox_simple_cpu0_to_cpu1_avmm_msg_sender.address
		.mailbox_simple_cpu0_to_cpu1_avmm_msg_sender_write             (mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_sender_write),          //                                                        .write
		.mailbox_simple_cpu0_to_cpu1_avmm_msg_sender_read              (mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_sender_read),           //                                                        .read
		.mailbox_simple_cpu0_to_cpu1_avmm_msg_sender_readdata          (mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_sender_readdata),       //                                                        .readdata
		.mailbox_simple_cpu0_to_cpu1_avmm_msg_sender_writedata         (mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_sender_writedata),      //                                                        .writedata
		.mailbox_simple_cpu0_to_cpu1_avmm_msg_sender_waitrequest       (mm_interconnect_0_mailbox_simple_cpu0_to_cpu1_avmm_msg_sender_waitrequest),    //                                                        .waitrequest
		.mailbox_simple_cpu1_to_cpu0_avmm_msg_receiver_address         (mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_receiver_address),      //           mailbox_simple_cpu1_to_cpu0_avmm_msg_receiver.address
		.mailbox_simple_cpu1_to_cpu0_avmm_msg_receiver_write           (mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_receiver_write),        //                                                        .write
		.mailbox_simple_cpu1_to_cpu0_avmm_msg_receiver_read            (mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_receiver_read),         //                                                        .read
		.mailbox_simple_cpu1_to_cpu0_avmm_msg_receiver_readdata        (mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_receiver_readdata),     //                                                        .readdata
		.mailbox_simple_cpu1_to_cpu0_avmm_msg_receiver_writedata       (mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_receiver_writedata),    //                                                        .writedata
		.mailbox_simple_cpu1_to_cpu0_avmm_msg_sender_address           (mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_sender_address),        //             mailbox_simple_cpu1_to_cpu0_avmm_msg_sender.address
		.mailbox_simple_cpu1_to_cpu0_avmm_msg_sender_write             (mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_sender_write),          //                                                        .write
		.mailbox_simple_cpu1_to_cpu0_avmm_msg_sender_read              (mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_sender_read),           //                                                        .read
		.mailbox_simple_cpu1_to_cpu0_avmm_msg_sender_readdata          (mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_sender_readdata),       //                                                        .readdata
		.mailbox_simple_cpu1_to_cpu0_avmm_msg_sender_writedata         (mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_sender_writedata),      //                                                        .writedata
		.mailbox_simple_cpu1_to_cpu0_avmm_msg_sender_waitrequest       (mm_interconnect_0_mailbox_simple_cpu1_to_cpu0_avmm_msg_sender_waitrequest),    //                                                        .waitrequest
		.mdma_from_idct_accel_csr_address                              (mm_interconnect_0_mdma_from_idct_accel_csr_address),                           //                                mdma_from_idct_accel_csr.address
		.mdma_from_idct_accel_csr_write                                (mm_interconnect_0_mdma_from_idct_accel_csr_write),                             //                                                        .write
		.mdma_from_idct_accel_csr_read                                 (mm_interconnect_0_mdma_from_idct_accel_csr_read),                              //                                                        .read
		.mdma_from_idct_accel_csr_readdata                             (mm_interconnect_0_mdma_from_idct_accel_csr_readdata),                          //                                                        .readdata
		.mdma_from_idct_accel_csr_writedata                            (mm_interconnect_0_mdma_from_idct_accel_csr_writedata),                         //                                                        .writedata
		.mdma_from_idct_accel_csr_byteenable                           (mm_interconnect_0_mdma_from_idct_accel_csr_byteenable),                        //                                                        .byteenable
		.mdma_from_idct_accel_descriptor_slave_write                   (mm_interconnect_0_mdma_from_idct_accel_descriptor_slave_write),                //                   mdma_from_idct_accel_descriptor_slave.write
		.mdma_from_idct_accel_descriptor_slave_writedata               (mm_interconnect_0_mdma_from_idct_accel_descriptor_slave_writedata),            //                                                        .writedata
		.mdma_from_idct_accel_descriptor_slave_byteenable              (mm_interconnect_0_mdma_from_idct_accel_descriptor_slave_byteenable),           //                                                        .byteenable
		.mdma_from_idct_accel_descriptor_slave_waitrequest             (mm_interconnect_0_mdma_from_idct_accel_descriptor_slave_waitrequest),          //                                                        .waitrequest
		.mdma_from_ycbcr_to_rgb_accel_csr_address                      (mm_interconnect_0_mdma_from_ycbcr_to_rgb_accel_csr_address),                   //                        mdma_from_ycbcr_to_rgb_accel_csr.address
		.mdma_from_ycbcr_to_rgb_accel_csr_write                        (mm_interconnect_0_mdma_from_ycbcr_to_rgb_accel_csr_write),                     //                                                        .write
		.mdma_from_ycbcr_to_rgb_accel_csr_read                         (mm_interconnect_0_mdma_from_ycbcr_to_rgb_accel_csr_read),                      //                                                        .read
		.mdma_from_ycbcr_to_rgb_accel_csr_readdata                     (mm_interconnect_0_mdma_from_ycbcr_to_rgb_accel_csr_readdata),                  //                                                        .readdata
		.mdma_from_ycbcr_to_rgb_accel_csr_writedata                    (mm_interconnect_0_mdma_from_ycbcr_to_rgb_accel_csr_writedata),                 //                                                        .writedata
		.mdma_from_ycbcr_to_rgb_accel_csr_byteenable                   (mm_interconnect_0_mdma_from_ycbcr_to_rgb_accel_csr_byteenable),                //                                                        .byteenable
		.mdma_from_ycbcr_to_rgb_accel_descriptor_slave_write           (mm_interconnect_0_mdma_from_ycbcr_to_rgb_accel_descriptor_slave_write),        //           mdma_from_ycbcr_to_rgb_accel_descriptor_slave.write
		.mdma_from_ycbcr_to_rgb_accel_descriptor_slave_writedata       (mm_interconnect_0_mdma_from_ycbcr_to_rgb_accel_descriptor_slave_writedata),    //                                                        .writedata
		.mdma_from_ycbcr_to_rgb_accel_descriptor_slave_byteenable      (mm_interconnect_0_mdma_from_ycbcr_to_rgb_accel_descriptor_slave_byteenable),   //                                                        .byteenable
		.mdma_from_ycbcr_to_rgb_accel_descriptor_slave_waitrequest     (mm_interconnect_0_mdma_from_ycbcr_to_rgb_accel_descriptor_slave_waitrequest),  //                                                        .waitrequest
		.mdma_to_idct_accel_csr_address                                (mm_interconnect_0_mdma_to_idct_accel_csr_address),                             //                                  mdma_to_idct_accel_csr.address
		.mdma_to_idct_accel_csr_write                                  (mm_interconnect_0_mdma_to_idct_accel_csr_write),                               //                                                        .write
		.mdma_to_idct_accel_csr_read                                   (mm_interconnect_0_mdma_to_idct_accel_csr_read),                                //                                                        .read
		.mdma_to_idct_accel_csr_readdata                               (mm_interconnect_0_mdma_to_idct_accel_csr_readdata),                            //                                                        .readdata
		.mdma_to_idct_accel_csr_writedata                              (mm_interconnect_0_mdma_to_idct_accel_csr_writedata),                           //                                                        .writedata
		.mdma_to_idct_accel_csr_byteenable                             (mm_interconnect_0_mdma_to_idct_accel_csr_byteenable),                          //                                                        .byteenable
		.mdma_to_idct_accel_descriptor_slave_write                     (mm_interconnect_0_mdma_to_idct_accel_descriptor_slave_write),                  //                     mdma_to_idct_accel_descriptor_slave.write
		.mdma_to_idct_accel_descriptor_slave_writedata                 (mm_interconnect_0_mdma_to_idct_accel_descriptor_slave_writedata),              //                                                        .writedata
		.mdma_to_idct_accel_descriptor_slave_byteenable                (mm_interconnect_0_mdma_to_idct_accel_descriptor_slave_byteenable),             //                                                        .byteenable
		.mdma_to_idct_accel_descriptor_slave_waitrequest               (mm_interconnect_0_mdma_to_idct_accel_descriptor_slave_waitrequest),            //                                                        .waitrequest
		.mdma_to_ycbcr_to_rgb_accel_cb_csr_address                     (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cb_csr_address),                  //                       mdma_to_ycbcr_to_rgb_accel_cb_csr.address
		.mdma_to_ycbcr_to_rgb_accel_cb_csr_write                       (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cb_csr_write),                    //                                                        .write
		.mdma_to_ycbcr_to_rgb_accel_cb_csr_read                        (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cb_csr_read),                     //                                                        .read
		.mdma_to_ycbcr_to_rgb_accel_cb_csr_readdata                    (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cb_csr_readdata),                 //                                                        .readdata
		.mdma_to_ycbcr_to_rgb_accel_cb_csr_writedata                   (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cb_csr_writedata),                //                                                        .writedata
		.mdma_to_ycbcr_to_rgb_accel_cb_csr_byteenable                  (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cb_csr_byteenable),               //                                                        .byteenable
		.mdma_to_ycbcr_to_rgb_accel_cb_descriptor_slave_write          (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cb_descriptor_slave_write),       //          mdma_to_ycbcr_to_rgb_accel_cb_descriptor_slave.write
		.mdma_to_ycbcr_to_rgb_accel_cb_descriptor_slave_writedata      (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cb_descriptor_slave_writedata),   //                                                        .writedata
		.mdma_to_ycbcr_to_rgb_accel_cb_descriptor_slave_byteenable     (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cb_descriptor_slave_byteenable),  //                                                        .byteenable
		.mdma_to_ycbcr_to_rgb_accel_cb_descriptor_slave_waitrequest    (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cb_descriptor_slave_waitrequest), //                                                        .waitrequest
		.mdma_to_ycbcr_to_rgb_accel_cr_csr_address                     (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cr_csr_address),                  //                       mdma_to_ycbcr_to_rgb_accel_cr_csr.address
		.mdma_to_ycbcr_to_rgb_accel_cr_csr_write                       (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cr_csr_write),                    //                                                        .write
		.mdma_to_ycbcr_to_rgb_accel_cr_csr_read                        (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cr_csr_read),                     //                                                        .read
		.mdma_to_ycbcr_to_rgb_accel_cr_csr_readdata                    (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cr_csr_readdata),                 //                                                        .readdata
		.mdma_to_ycbcr_to_rgb_accel_cr_csr_writedata                   (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cr_csr_writedata),                //                                                        .writedata
		.mdma_to_ycbcr_to_rgb_accel_cr_csr_byteenable                  (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cr_csr_byteenable),               //                                                        .byteenable
		.mdma_to_ycbcr_to_rgb_accel_cr_descriptor_slave_write          (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cr_descriptor_slave_write),       //          mdma_to_ycbcr_to_rgb_accel_cr_descriptor_slave.write
		.mdma_to_ycbcr_to_rgb_accel_cr_descriptor_slave_writedata      (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cr_descriptor_slave_writedata),   //                                                        .writedata
		.mdma_to_ycbcr_to_rgb_accel_cr_descriptor_slave_byteenable     (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cr_descriptor_slave_byteenable),  //                                                        .byteenable
		.mdma_to_ycbcr_to_rgb_accel_cr_descriptor_slave_waitrequest    (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_cr_descriptor_slave_waitrequest), //                                                        .waitrequest
		.mdma_to_ycbcr_to_rgb_accel_y_csr_address                      (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_y_csr_address),                   //                        mdma_to_ycbcr_to_rgb_accel_y_csr.address
		.mdma_to_ycbcr_to_rgb_accel_y_csr_write                        (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_y_csr_write),                     //                                                        .write
		.mdma_to_ycbcr_to_rgb_accel_y_csr_read                         (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_y_csr_read),                      //                                                        .read
		.mdma_to_ycbcr_to_rgb_accel_y_csr_readdata                     (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_y_csr_readdata),                  //                                                        .readdata
		.mdma_to_ycbcr_to_rgb_accel_y_csr_writedata                    (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_y_csr_writedata),                 //                                                        .writedata
		.mdma_to_ycbcr_to_rgb_accel_y_csr_byteenable                   (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_y_csr_byteenable),                //                                                        .byteenable
		.mdma_to_ycbcr_to_rgb_accel_y_descriptor_slave_write           (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_y_descriptor_slave_write),        //           mdma_to_ycbcr_to_rgb_accel_y_descriptor_slave.write
		.mdma_to_ycbcr_to_rgb_accel_y_descriptor_slave_writedata       (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_y_descriptor_slave_writedata),    //                                                        .writedata
		.mdma_to_ycbcr_to_rgb_accel_y_descriptor_slave_byteenable      (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_y_descriptor_slave_byteenable),   //                                                        .byteenable
		.mdma_to_ycbcr_to_rgb_accel_y_descriptor_slave_waitrequest     (mm_interconnect_0_mdma_to_ycbcr_to_rgb_accel_y_descriptor_slave_waitrequest),  //                                                        .waitrequest
		.mutex_0_s1_address                                            (mm_interconnect_0_mutex_0_s1_address),                                         //                                              mutex_0_s1.address
		.mutex_0_s1_write                                              (mm_interconnect_0_mutex_0_s1_write),                                           //                                                        .write
		.mutex_0_s1_read                                               (mm_interconnect_0_mutex_0_s1_read),                                            //                                                        .read
		.mutex_0_s1_readdata                                           (mm_interconnect_0_mutex_0_s1_readdata),                                        //                                                        .readdata
		.mutex_0_s1_writedata                                          (mm_interconnect_0_mutex_0_s1_writedata),                                       //                                                        .writedata
		.mutex_0_s1_chipselect                                         (mm_interconnect_0_mutex_0_s1_chipselect),                                      //                                                        .chipselect
		.sd_cont_slave_address                                         (mm_interconnect_0_sd_cont_slave_address),                                      //                                           sd_cont_slave.address
		.sd_cont_slave_write                                           (mm_interconnect_0_sd_cont_slave_write),                                        //                                                        .write
		.sd_cont_slave_read                                            (mm_interconnect_0_sd_cont_slave_read),                                         //                                                        .read
		.sd_cont_slave_readdata                                        (mm_interconnect_0_sd_cont_slave_readdata),                                     //                                                        .readdata
		.sd_cont_slave_writedata                                       (mm_interconnect_0_sd_cont_slave_writedata),                                    //                                                        .writedata
		.sd_cont_slave_waitrequest                                     (~mm_interconnect_0_sd_cont_slave_waitrequest),                                 //                                                        .waitrequest
		.sd_cont_slave_chipselect                                      (mm_interconnect_0_sd_cont_slave_chipselect),                                   //                                                        .chipselect
		.sram_uas_address                                              (mm_interconnect_0_sram_uas_address),                                           //                                                sram_uas.address
		.sram_uas_write                                                (mm_interconnect_0_sram_uas_write),                                             //                                                        .write
		.sram_uas_read                                                 (mm_interconnect_0_sram_uas_read),                                              //                                                        .read
		.sram_uas_readdata                                             (mm_interconnect_0_sram_uas_readdata),                                          //                                                        .readdata
		.sram_uas_writedata                                            (mm_interconnect_0_sram_uas_writedata),                                         //                                                        .writedata
		.sram_uas_burstcount                                           (mm_interconnect_0_sram_uas_burstcount),                                        //                                                        .burstcount
		.sram_uas_byteenable                                           (mm_interconnect_0_sram_uas_byteenable),                                        //                                                        .byteenable
		.sram_uas_readdatavalid                                        (mm_interconnect_0_sram_uas_readdatavalid),                                     //                                                        .readdatavalid
		.sram_uas_waitrequest                                          (mm_interconnect_0_sram_uas_waitrequest),                                       //                                                        .waitrequest
		.sram_uas_lock                                                 (mm_interconnect_0_sram_uas_lock),                                              //                                                        .lock
		.sram_uas_debugaccess                                          (mm_interconnect_0_sram_uas_debugaccess),                                       //                                                        .debugaccess
		.sysid_control_slave_address                                   (mm_interconnect_0_sysid_control_slave_address),                                //                                     sysid_control_slave.address
		.sysid_control_slave_readdata                                  (mm_interconnect_0_sysid_control_slave_readdata),                               //                                                        .readdata
		.timer_0_0_s1_address                                          (mm_interconnect_0_timer_0_0_s1_address),                                       //                                            timer_0_0_s1.address
		.timer_0_0_s1_write                                            (mm_interconnect_0_timer_0_0_s1_write),                                         //                                                        .write
		.timer_0_0_s1_readdata                                         (mm_interconnect_0_timer_0_0_s1_readdata),                                      //                                                        .readdata
		.timer_0_0_s1_writedata                                        (mm_interconnect_0_timer_0_0_s1_writedata),                                     //                                                        .writedata
		.timer_0_0_s1_chipselect                                       (mm_interconnect_0_timer_0_0_s1_chipselect),                                    //                                                        .chipselect
		.timer_0_1_s1_address                                          (mm_interconnect_0_timer_0_1_s1_address),                                       //                                            timer_0_1_s1.address
		.timer_0_1_s1_write                                            (mm_interconnect_0_timer_0_1_s1_write),                                         //                                                        .write
		.timer_0_1_s1_readdata                                         (mm_interconnect_0_timer_0_1_s1_readdata),                                      //                                                        .readdata
		.timer_0_1_s1_writedata                                        (mm_interconnect_0_timer_0_1_s1_writedata),                                     //                                                        .writedata
		.timer_0_1_s1_chipselect                                       (mm_interconnect_0_timer_0_1_s1_chipselect),                                    //                                                        .chipselect
		.timer_1_0_s1_address                                          (mm_interconnect_0_timer_1_0_s1_address),                                       //                                            timer_1_0_s1.address
		.timer_1_0_s1_write                                            (mm_interconnect_0_timer_1_0_s1_write),                                         //                                                        .write
		.timer_1_0_s1_readdata                                         (mm_interconnect_0_timer_1_0_s1_readdata),                                      //                                                        .readdata
		.timer_1_0_s1_writedata                                        (mm_interconnect_0_timer_1_0_s1_writedata),                                     //                                                        .writedata
		.timer_1_0_s1_chipselect                                       (mm_interconnect_0_timer_1_0_s1_chipselect),                                    //                                                        .chipselect
		.timer_1_1_s1_address                                          (mm_interconnect_0_timer_1_1_s1_address),                                       //                                            timer_1_1_s1.address
		.timer_1_1_s1_write                                            (mm_interconnect_0_timer_1_1_s1_write),                                         //                                                        .write
		.timer_1_1_s1_readdata                                         (mm_interconnect_0_timer_1_1_s1_readdata),                                      //                                                        .readdata
		.timer_1_1_s1_writedata                                        (mm_interconnect_0_timer_1_1_s1_writedata),                                     //                                                        .writedata
		.timer_1_1_s1_chipselect                                       (mm_interconnect_0_timer_1_1_s1_chipselect),                                    //                                                        .chipselect
		.video_dma_csr_address                                         (mm_interconnect_0_video_dma_csr_address),                                      //                                           video_dma_csr.address
		.video_dma_csr_write                                           (mm_interconnect_0_video_dma_csr_write),                                        //                                                        .write
		.video_dma_csr_read                                            (mm_interconnect_0_video_dma_csr_read),                                         //                                                        .read
		.video_dma_csr_readdata                                        (mm_interconnect_0_video_dma_csr_readdata),                                     //                                                        .readdata
		.video_dma_csr_writedata                                       (mm_interconnect_0_video_dma_csr_writedata),                                    //                                                        .writedata
		.video_dma_csr_byteenable                                      (mm_interconnect_0_video_dma_csr_byteenable),                                   //                                                        .byteenable
		.video_dma_descriptor_slave_write                              (mm_interconnect_0_video_dma_descriptor_slave_write),                           //                              video_dma_descriptor_slave.write
		.video_dma_descriptor_slave_writedata                          (mm_interconnect_0_video_dma_descriptor_slave_writedata),                       //                                                        .writedata
		.video_dma_descriptor_slave_byteenable                         (mm_interconnect_0_video_dma_descriptor_slave_byteenable),                      //                                                        .byteenable
		.video_dma_descriptor_slave_waitrequest                        (mm_interconnect_0_video_dma_descriptor_slave_waitrequest)                      //                                                        .waitrequest
	);

	ECE423_QSYS_mm_interconnect_1 mm_interconnect_1 (
		.clk_125_clk_clk                                     (clk_125_clk),                                         //                                   clk_125_clk.clk
		.lpddr2_mp_cmd_reset_n_1_reset_bridge_in_reset_reset (reset_controller_0_reset_out_reset),                  // lpddr2_mp_cmd_reset_n_1_reset_bridge_in_reset.reset
		.video_dma_reset_n_reset_bridge_in_reset_reset       (reset_controller_0_reset_out_reset),                  //       video_dma_reset_n_reset_bridge_in_reset.reset
		.mdma_to_idct_accel_mm_read_address                  (mdma_to_idct_accel_mm_read_address),                  //                    mdma_to_idct_accel_mm_read.address
		.mdma_to_idct_accel_mm_read_waitrequest              (mdma_to_idct_accel_mm_read_waitrequest),              //                                              .waitrequest
		.mdma_to_idct_accel_mm_read_burstcount               (mdma_to_idct_accel_mm_read_burstcount),               //                                              .burstcount
		.mdma_to_idct_accel_mm_read_byteenable               (mdma_to_idct_accel_mm_read_byteenable),               //                                              .byteenable
		.mdma_to_idct_accel_mm_read_read                     (mdma_to_idct_accel_mm_read_read),                     //                                              .read
		.mdma_to_idct_accel_mm_read_readdata                 (mdma_to_idct_accel_mm_read_readdata),                 //                                              .readdata
		.mdma_to_idct_accel_mm_read_readdatavalid            (mdma_to_idct_accel_mm_read_readdatavalid),            //                                              .readdatavalid
		.mdma_to_ycbcr_to_rgb_accel_cb_mm_read_address       (mdma_to_ycbcr_to_rgb_accel_cb_mm_read_address),       //         mdma_to_ycbcr_to_rgb_accel_cb_mm_read.address
		.mdma_to_ycbcr_to_rgb_accel_cb_mm_read_waitrequest   (mdma_to_ycbcr_to_rgb_accel_cb_mm_read_waitrequest),   //                                              .waitrequest
		.mdma_to_ycbcr_to_rgb_accel_cb_mm_read_burstcount    (mdma_to_ycbcr_to_rgb_accel_cb_mm_read_burstcount),    //                                              .burstcount
		.mdma_to_ycbcr_to_rgb_accel_cb_mm_read_byteenable    (mdma_to_ycbcr_to_rgb_accel_cb_mm_read_byteenable),    //                                              .byteenable
		.mdma_to_ycbcr_to_rgb_accel_cb_mm_read_read          (mdma_to_ycbcr_to_rgb_accel_cb_mm_read_read),          //                                              .read
		.mdma_to_ycbcr_to_rgb_accel_cb_mm_read_readdata      (mdma_to_ycbcr_to_rgb_accel_cb_mm_read_readdata),      //                                              .readdata
		.mdma_to_ycbcr_to_rgb_accel_cb_mm_read_readdatavalid (mdma_to_ycbcr_to_rgb_accel_cb_mm_read_readdatavalid), //                                              .readdatavalid
		.mdma_to_ycbcr_to_rgb_accel_cr_mm_read_address       (mdma_to_ycbcr_to_rgb_accel_cr_mm_read_address),       //         mdma_to_ycbcr_to_rgb_accel_cr_mm_read.address
		.mdma_to_ycbcr_to_rgb_accel_cr_mm_read_waitrequest   (mdma_to_ycbcr_to_rgb_accel_cr_mm_read_waitrequest),   //                                              .waitrequest
		.mdma_to_ycbcr_to_rgb_accel_cr_mm_read_burstcount    (mdma_to_ycbcr_to_rgb_accel_cr_mm_read_burstcount),    //                                              .burstcount
		.mdma_to_ycbcr_to_rgb_accel_cr_mm_read_byteenable    (mdma_to_ycbcr_to_rgb_accel_cr_mm_read_byteenable),    //                                              .byteenable
		.mdma_to_ycbcr_to_rgb_accel_cr_mm_read_read          (mdma_to_ycbcr_to_rgb_accel_cr_mm_read_read),          //                                              .read
		.mdma_to_ycbcr_to_rgb_accel_cr_mm_read_readdata      (mdma_to_ycbcr_to_rgb_accel_cr_mm_read_readdata),      //                                              .readdata
		.mdma_to_ycbcr_to_rgb_accel_cr_mm_read_readdatavalid (mdma_to_ycbcr_to_rgb_accel_cr_mm_read_readdatavalid), //                                              .readdatavalid
		.mdma_to_ycbcr_to_rgb_accel_y_mm_read_address        (mdma_to_ycbcr_to_rgb_accel_y_mm_read_address),        //          mdma_to_ycbcr_to_rgb_accel_y_mm_read.address
		.mdma_to_ycbcr_to_rgb_accel_y_mm_read_waitrequest    (mdma_to_ycbcr_to_rgb_accel_y_mm_read_waitrequest),    //                                              .waitrequest
		.mdma_to_ycbcr_to_rgb_accel_y_mm_read_burstcount     (mdma_to_ycbcr_to_rgb_accel_y_mm_read_burstcount),     //                                              .burstcount
		.mdma_to_ycbcr_to_rgb_accel_y_mm_read_byteenable     (mdma_to_ycbcr_to_rgb_accel_y_mm_read_byteenable),     //                                              .byteenable
		.mdma_to_ycbcr_to_rgb_accel_y_mm_read_read           (mdma_to_ycbcr_to_rgb_accel_y_mm_read_read),           //                                              .read
		.mdma_to_ycbcr_to_rgb_accel_y_mm_read_readdata       (mdma_to_ycbcr_to_rgb_accel_y_mm_read_readdata),       //                                              .readdata
		.mdma_to_ycbcr_to_rgb_accel_y_mm_read_readdatavalid  (mdma_to_ycbcr_to_rgb_accel_y_mm_read_readdatavalid),  //                                              .readdatavalid
		.video_dma_mm_read_address                           (video_dma_mm_read_address),                           //                             video_dma_mm_read.address
		.video_dma_mm_read_waitrequest                       (video_dma_mm_read_waitrequest),                       //                                              .waitrequest
		.video_dma_mm_read_burstcount                        (video_dma_mm_read_burstcount),                        //                                              .burstcount
		.video_dma_mm_read_byteenable                        (video_dma_mm_read_byteenable),                        //                                              .byteenable
		.video_dma_mm_read_read                              (video_dma_mm_read_read),                              //                                              .read
		.video_dma_mm_read_readdata                          (video_dma_mm_read_readdata),                          //                                              .readdata
		.video_dma_mm_read_readdatavalid                     (video_dma_mm_read_readdatavalid),                     //                                              .readdatavalid
		.lpddr2_avl_1_address                                (mm_interconnect_1_lpddr2_avl_1_address),              //                                  lpddr2_avl_1.address
		.lpddr2_avl_1_write                                  (mm_interconnect_1_lpddr2_avl_1_write),                //                                              .write
		.lpddr2_avl_1_read                                   (mm_interconnect_1_lpddr2_avl_1_read),                 //                                              .read
		.lpddr2_avl_1_readdata                               (mm_interconnect_1_lpddr2_avl_1_readdata),             //                                              .readdata
		.lpddr2_avl_1_writedata                              (mm_interconnect_1_lpddr2_avl_1_writedata),            //                                              .writedata
		.lpddr2_avl_1_beginbursttransfer                     (mm_interconnect_1_lpddr2_avl_1_beginbursttransfer),   //                                              .beginbursttransfer
		.lpddr2_avl_1_burstcount                             (mm_interconnect_1_lpddr2_avl_1_burstcount),           //                                              .burstcount
		.lpddr2_avl_1_byteenable                             (mm_interconnect_1_lpddr2_avl_1_byteenable),           //                                              .byteenable
		.lpddr2_avl_1_readdatavalid                          (mm_interconnect_1_lpddr2_avl_1_readdatavalid),        //                                              .readdatavalid
		.lpddr2_avl_1_waitrequest                            (~mm_interconnect_1_lpddr2_avl_1_waitrequest)          //                                              .waitrequest
	);

	ECE423_QSYS_mm_interconnect_2 mm_interconnect_2 (
		.clk_125_clk_clk                                          (clk_125_clk),                                       //                                        clk_125_clk.clk
		.lpddr2_mp_cmd_reset_n_2_reset_bridge_in_reset_reset      (reset_controller_0_reset_out_reset),                //      lpddr2_mp_cmd_reset_n_2_reset_bridge_in_reset.reset
		.mdma_from_idct_accel_reset_n_reset_bridge_in_reset_reset (reset_controller_0_reset_out_reset),                // mdma_from_idct_accel_reset_n_reset_bridge_in_reset.reset
		.mdma_from_idct_accel_mm_write_address                    (mdma_from_idct_accel_mm_write_address),             //                      mdma_from_idct_accel_mm_write.address
		.mdma_from_idct_accel_mm_write_waitrequest                (mdma_from_idct_accel_mm_write_waitrequest),         //                                                   .waitrequest
		.mdma_from_idct_accel_mm_write_burstcount                 (mdma_from_idct_accel_mm_write_burstcount),          //                                                   .burstcount
		.mdma_from_idct_accel_mm_write_byteenable                 (mdma_from_idct_accel_mm_write_byteenable),          //                                                   .byteenable
		.mdma_from_idct_accel_mm_write_write                      (mdma_from_idct_accel_mm_write_write),               //                                                   .write
		.mdma_from_idct_accel_mm_write_writedata                  (mdma_from_idct_accel_mm_write_writedata),           //                                                   .writedata
		.mdma_from_ycbcr_to_rgb_accel_mm_write_address            (mdma_from_ycbcr_to_rgb_accel_mm_write_address),     //              mdma_from_ycbcr_to_rgb_accel_mm_write.address
		.mdma_from_ycbcr_to_rgb_accel_mm_write_waitrequest        (mdma_from_ycbcr_to_rgb_accel_mm_write_waitrequest), //                                                   .waitrequest
		.mdma_from_ycbcr_to_rgb_accel_mm_write_burstcount         (mdma_from_ycbcr_to_rgb_accel_mm_write_burstcount),  //                                                   .burstcount
		.mdma_from_ycbcr_to_rgb_accel_mm_write_byteenable         (mdma_from_ycbcr_to_rgb_accel_mm_write_byteenable),  //                                                   .byteenable
		.mdma_from_ycbcr_to_rgb_accel_mm_write_write              (mdma_from_ycbcr_to_rgb_accel_mm_write_write),       //                                                   .write
		.mdma_from_ycbcr_to_rgb_accel_mm_write_writedata          (mdma_from_ycbcr_to_rgb_accel_mm_write_writedata),   //                                                   .writedata
		.lpddr2_avl_2_address                                     (mm_interconnect_2_lpddr2_avl_2_address),            //                                       lpddr2_avl_2.address
		.lpddr2_avl_2_write                                       (mm_interconnect_2_lpddr2_avl_2_write),              //                                                   .write
		.lpddr2_avl_2_read                                        (mm_interconnect_2_lpddr2_avl_2_read),               //                                                   .read
		.lpddr2_avl_2_readdata                                    (mm_interconnect_2_lpddr2_avl_2_readdata),           //                                                   .readdata
		.lpddr2_avl_2_writedata                                   (mm_interconnect_2_lpddr2_avl_2_writedata),          //                                                   .writedata
		.lpddr2_avl_2_beginbursttransfer                          (mm_interconnect_2_lpddr2_avl_2_beginbursttransfer), //                                                   .beginbursttransfer
		.lpddr2_avl_2_burstcount                                  (mm_interconnect_2_lpddr2_avl_2_burstcount),         //                                                   .burstcount
		.lpddr2_avl_2_byteenable                                  (mm_interconnect_2_lpddr2_avl_2_byteenable),         //                                                   .byteenable
		.lpddr2_avl_2_readdatavalid                               (mm_interconnect_2_lpddr2_avl_2_readdatavalid),      //                                                   .readdatavalid
		.lpddr2_avl_2_waitrequest                                 (~mm_interconnect_2_lpddr2_avl_2_waitrequest)        //                                                   .waitrequest
	);

	ECE423_QSYS_irq_mapper irq_mapper (
		.clk           (clk_125_clk),                    //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),       // receiver6.irq
		.sender_irq    (cpu_0_irq_irq)                   //    sender.irq
	);

	ECE423_QSYS_irq_mapper_001 irq_mapper_001 (
		.clk            (clk_125_clk),                        //        clk.clk
		.reset          (rst_controller_001_reset_out_reset), //  clk_reset.reset
		.receiver0_irq  (irq_mapper_001_receiver0_irq),       //  receiver0.irq
		.receiver1_irq  (irq_mapper_001_receiver1_irq),       //  receiver1.irq
		.receiver2_irq  (irq_mapper_001_receiver2_irq),       //  receiver2.irq
		.receiver3_irq  (irq_mapper_001_receiver3_irq),       //  receiver3.irq
		.receiver4_irq  (irq_mapper_001_receiver4_irq),       //  receiver4.irq
		.receiver5_irq  (irq_mapper_001_receiver5_irq),       //  receiver5.irq
		.receiver6_irq  (irq_mapper_001_receiver6_irq),       //  receiver6.irq
		.receiver7_irq  (irq_mapper_001_receiver7_irq),       //  receiver7.irq
		.receiver8_irq  (irq_mapper_001_receiver8_irq),       //  receiver8.irq
		.receiver9_irq  (irq_mapper_001_receiver9_irq),       //  receiver9.irq
		.receiver10_irq (irq_mapper_001_receiver10_irq),      // receiver10.irq
		.sender_irq     (cpu_1_irq_irq)                       //     sender.irq
	);

	ECE423_QSYS_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (1),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (video_clk_clk),                         // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_002_reset_out_reset),    // in_rst_0.reset
		.in_0_data           (video_fifo_out_data),                   //     in_0.data
		.in_0_valid          (video_fifo_out_valid),                  //         .valid
		.in_0_ready          (video_fifo_out_ready),                  //         .ready
		.in_0_startofpacket  (video_fifo_out_startofpacket),          //         .startofpacket
		.in_0_endofpacket    (video_fifo_out_endofpacket),            //         .endofpacket
		.in_0_empty          (video_fifo_out_empty),                  //         .empty
		.out_0_data          (avalon_st_adapter_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_out_0_empty)          //         .empty
	);

	ECE423_QSYS_avalon_st_adapter_001 #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (1)
	) avalon_st_adapter_001 (
		.in_clk_0_clk        (clk_125_clk),                               // in_clk_0.clk
		.in_rst_0_reset      (reset_controller_0_reset_out_reset),        // in_rst_0.reset
		.in_0_data           (video_dma_st_source_data),                  //     in_0.data
		.in_0_valid          (video_dma_st_source_valid),                 //         .valid
		.in_0_ready          (video_dma_st_source_ready),                 //         .ready
		.in_0_startofpacket  (video_dma_st_source_startofpacket),         //         .startofpacket
		.in_0_endofpacket    (video_dma_st_source_endofpacket),           //         .endofpacket
		.in_0_empty          (video_dma_st_source_empty),                 //         .empty
		.out_0_data          (avalon_st_adapter_001_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_001_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_001_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_001_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_001_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_001_out_0_empty)          //         .empty
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (cpu_0_debug_reset_request_reset),    // reset_in0.reset
		.reset_in1      (reset_controller_0_reset_out_reset), // reset_in1.reset
		.clk            (clk_125_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (cpu_1_debug_reset_request_reset),        // reset_in0.reset
		.reset_in1      (reset_controller_0_reset_out_reset),     // reset_in1.reset
		.clk            (clk_125_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (reset_controller_0_reset_out_reset), // reset_in0.reset
		.clk            (video_clk_clk),                      //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (reset_controller_0_reset_out_reset), // reset_in0.reset
		.clk            (clk_50_clk),                         //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
